`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:54:50 01/19/2015 
// Design Name: 
// Module Name:    rand_table_7 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module rand_table_9(axi_aclk , axi_aresetn , index_num , rand_out , en);
	input			axi_aclk , axi_aresetn , en;
	input		[7:0]	index_num;
	output		[31:0]	rand_out;

	reg 		[31:0]	random_num_table  [255:0];

	assign rand_out = en?random_num_table[index_num]:32'd0;
	
	always@(posedge axi_aclk)
	begin
		random_num_table[0]  <= 32'b	00001001011011001000010010000110	;
		random_num_table[1]  <= 32'b	00001010111010101010101110000011	;
		random_num_table[2]  <= 32'b	00011011001001101000111010100011	;
		random_num_table[3]  <= 32'b	00000101110000010001100101101000	;
		random_num_table[4]  <= 32'b	00001000010100110011010011000010	;
		random_num_table[5]  <= 32'b	00000000100011111111001001101100	;
		random_num_table[6]  <= 32'b	00010111000010111001100001001101	;
		random_num_table[7]  <= 32'b	00001001010101111000100010010000	;
		random_num_table[8]  <= 32'b	00011101010010000011001100011011	;
		random_num_table[9]  <= 32'b	00010110100111001101001010100001	;
		random_num_table[10]  <= 32'b	00010101110001110100000000000000	;
		random_num_table[11]  <= 32'b	00011011101100000010111110100001	;
		random_num_table[12]  <= 32'b	00011100100010011001110011101010	;
		random_num_table[13]  <= 32'b	00010101011111001100111001010100	;
		random_num_table[14]  <= 32'b	00000000011001000101110010010000	;
		random_num_table[15]  <= 32'b	00000100101011100101111111110001	;
		random_num_table[16]  <= 32'b	00010110010010001100101110000000	;
		random_num_table[17]  <= 32'b	00000001110011111111111010000100	;
		random_num_table[18]  <= 32'b	00001111101100111110110010010011	;
		random_num_table[19]  <= 32'b	00000110001000110111111010101100	;
		random_num_table[20]  <= 32'b	00010001111101111000101111111010	;
		random_num_table[21]  <= 32'b	00011111100101011111100110100000	;
		random_num_table[22]  <= 32'b	00000110011111011100010100101101	;
		random_num_table[23]  <= 32'b	00011100001001100011001110000101	;
		random_num_table[24]  <= 32'b	00011001001111000101010110011111	;
		random_num_table[25]  <= 32'b	00001000011100111010001000100101	;
		random_num_table[26]  <= 32'b	00010011101100011111011011100111	;
		random_num_table[27]  <= 32'b	00000110010000001011111100001001	;
		random_num_table[28]  <= 32'b	00000001110111110011010111000101	;
		random_num_table[29]  <= 32'b	00011100111000001111001011101000	;
		random_num_table[30]  <= 32'b	00010101000111000011001010100111	;
		random_num_table[31]  <= 32'b	00011111001011010110000010001110	;
		random_num_table[32]  <= 32'b	00000101011011000001010110110110	;
		random_num_table[33]  <= 32'b	00010000101001011000010011011010	;
		random_num_table[34]  <= 32'b	00011010101011001110101110100000	;
		random_num_table[35]  <= 32'b	00000101111110010011101110001000	;
		random_num_table[36]  <= 32'b	00010110000001011100111110000100	;
		random_num_table[37]  <= 32'b	00011110111101100110011000100101	;
		random_num_table[38]  <= 32'b	00010101111111101111100001000111	;
		random_num_table[39]  <= 32'b	00001101001101001011111100000000	;
		random_num_table[40]  <= 32'b	00001110011110111110010000110001	;
		random_num_table[41]  <= 32'b	00001000010101110000010111110111	;
		random_num_table[42]  <= 32'b	00001101001110001011010001100001	;
		random_num_table[43]  <= 32'b	00001111100010100111001010010001	;
		random_num_table[44]  <= 32'b	00000000111100001110110010111101	;
		random_num_table[45]  <= 32'b	00000011011100010110100001101011	;
		random_num_table[46]  <= 32'b	00011101101010011010010010101001	;
		random_num_table[47]  <= 32'b	00001101101011001000010110010001	;
		random_num_table[48]  <= 32'b	00001110110100100010111010111111	;
		random_num_table[49]  <= 32'b	00011010001010110001111101000000	;
		random_num_table[50]  <= 32'b	00010111001001110010010100010000	;
		random_num_table[51]  <= 32'b	00011110011011011100011011101101	;
		random_num_table[52]  <= 32'b	00000111010111110001000100000110	;
		random_num_table[53]  <= 32'b	00001100011100011011111000101010	;
		random_num_table[54]  <= 32'b	00011011100010000111110100110101	;
		random_num_table[55]  <= 32'b	00001000001010101001100010001110	;
		random_num_table[56]  <= 32'b	00010000100001111000101011100100	;
		random_num_table[57]  <= 32'b	00000110101110000110000001000001	;
		random_num_table[58]  <= 32'b	00011100011011011011111010111110	;
		random_num_table[59]  <= 32'b	00001111010010110000000001001001	;
		random_num_table[60]  <= 32'b	00000101000000100001111000111110	;
		random_num_table[61]  <= 32'b	00011001111001111000110110110110	;
		random_num_table[62]  <= 32'b	00001101100101101001000000011010	;
		random_num_table[63]  <= 32'b	00011111100100110110011000011111	;
		random_num_table[64]  <= 32'b	00000101111000111111101011011011	;
		random_num_table[65]  <= 32'b	00001001100010110110001100100010	;
		random_num_table[66]  <= 32'b	00000111010001111000000011010111	;
		random_num_table[67]  <= 32'b	00011100111001001011100010001101	;
		random_num_table[68]  <= 32'b	00000000100000001101000001101011	;
		random_num_table[69]  <= 32'b	00010100110011001010110101111000	;
		random_num_table[70]  <= 32'b	00010000011111111011100000101011	;
		random_num_table[71]  <= 32'b	00011011110010010101110100100000	;
		random_num_table[72]  <= 32'b	00001100101101011000110111100001	;
		random_num_table[73]  <= 32'b	00001011011101010110111100111100	;
		random_num_table[74]  <= 32'b	00011101010100001101110111111000	;
		random_num_table[75]  <= 32'b	00011101011101111100010010001100	;
		random_num_table[76]  <= 32'b	00000000100111100111010000100101	;
		random_num_table[77]  <= 32'b	00010110111001101010100100100100	;
		random_num_table[78]  <= 32'b	00000011001001011100001011101101	;
		random_num_table[79]  <= 32'b	00010101010010000000111101100011	;
		random_num_table[80]  <= 32'b	00001001010100110011011011110100	;
		random_num_table[81]  <= 32'b	00001111000010000110000001010100	;
		random_num_table[82]  <= 32'b	00011001101111111001011011001111	;
		random_num_table[83]  <= 32'b	00001111000101011110010101110001	;
		random_num_table[84]  <= 32'b	00011000001100010101011000110111	;
		random_num_table[85]  <= 32'b	00010100111000100110111101100011	;
		random_num_table[86]  <= 32'b	00010001010000111101110011101000	;
		random_num_table[87]  <= 32'b	00001011001001110000101011011101	;
		random_num_table[88]  <= 32'b	00001101000010011110000100101110	;
		random_num_table[89]  <= 32'b	00010111000101001001100010010110	;
		random_num_table[90]  <= 32'b	00000001110011010010110111111001	;
		random_num_table[91]  <= 32'b	00000000010000001000011111100111	;
		random_num_table[92]  <= 32'b	00011100101011110011000110011011	;
		random_num_table[93]  <= 32'b	00011000100010101111111110000110	;
		random_num_table[94]  <= 32'b	00000101100101101000100001100001	;
		random_num_table[95]  <= 32'b	00011111110000101001111001010010	;
		random_num_table[96]  <= 32'b	00011001110011000001101101110111	;
		random_num_table[97]  <= 32'b	00001010000001000111000011001111	;
		random_num_table[98]  <= 32'b	00011000110000000000000101101000	;
		random_num_table[99]  <= 32'b	00000111010110101000001110000100	;
		random_num_table[100]  <= 32'b	00010011000111001100000000001011	;
		random_num_table[101]  <= 32'b	00010000111101101010100111010101	;
		random_num_table[102]  <= 32'b	00000001000010011000110000001111	;
		random_num_table[103]  <= 32'b	00001101000100100100100110001110	;
		random_num_table[104]  <= 32'b	00011000110011000101100000000001	;
		random_num_table[105]  <= 32'b	00011010000100111010000011010010	;
		random_num_table[106]  <= 32'b	00000111101011111011101001001001	;
		random_num_table[107]  <= 32'b	00001100110000001001011011100001	;
		random_num_table[108]  <= 32'b	00010001100111100100001100010110	;
		random_num_table[109]  <= 32'b	00001000101001100101001100100101	;
		random_num_table[110]  <= 32'b	00000010110001010100001110011000	;
		random_num_table[111]  <= 32'b	00000110111111100010001111100010	;
		random_num_table[112]  <= 32'b	00001101010101111110110011010101	;
		random_num_table[113]  <= 32'b	00001011011010011110101111111101	;
		random_num_table[114]  <= 32'b	00010100111100010011110111101000	;
		random_num_table[115]  <= 32'b	00010111011110000111100011011101	;
		random_num_table[116]  <= 32'b	00011001111111101010100000001000	;
		random_num_table[117]  <= 32'b	00011011101100011001000110000000	;
		random_num_table[118]  <= 32'b	00011000101100110011010111111010	;
		random_num_table[119]  <= 32'b	00001100000111001000101101101110	;
		random_num_table[120]  <= 32'b	00011100111111111001001110101100	;
		random_num_table[121]  <= 32'b	00011111001111100101101100101100	;
		random_num_table[122]  <= 32'b	00010101010110001001110011100111	;
		random_num_table[123]  <= 32'b	00001100100111100001000010111111	;
		random_num_table[124]  <= 32'b	00011101111000000101011110101001	;
		random_num_table[125]  <= 32'b	00000100100011011011110101011010	;
		random_num_table[126]  <= 32'b	00010110001100000111111000100110	;
		random_num_table[127]  <= 32'b	00011100110010100101100001101010	;
		random_num_table[128]  <= 32'b	00000000010110011101010000011000	;
		random_num_table[129]  <= 32'b	00011001101100001100000000001110	;
		random_num_table[130]  <= 32'b	00000111100110111101110101100100	;
		random_num_table[131]  <= 32'b	00011001111110000111111111110001	;
		random_num_table[132]  <= 32'b	00001010101001111010110001101110	;
		random_num_table[133]  <= 32'b	00000101010001010101001011010101	;
		random_num_table[134]  <= 32'b	00010001110000001011001000100110	;
		random_num_table[135]  <= 32'b	00001011111101011110100101100110	;
		random_num_table[136]  <= 32'b	00001110110111100111101111011110	;
		random_num_table[137]  <= 32'b	00010010011110011010110100000010	;
		random_num_table[138]  <= 32'b	00001001011000100110001111010001	;
		random_num_table[139]  <= 32'b	00010110011100011010111100011011	;
		random_num_table[140]  <= 32'b	00010111010100100110010111010001	;
		random_num_table[141]  <= 32'b	00001001000010101011000100111011	;
		random_num_table[142]  <= 32'b	00001001011000100101000001011010	;
		random_num_table[143]  <= 32'b	00000100100011101101110100110001	;
		random_num_table[144]  <= 32'b	00010110111010101111000011100110	;
		random_num_table[145]  <= 32'b	00010000100010111111100100001111	;
		random_num_table[146]  <= 32'b	00000000011000010110101110010101	;
		random_num_table[147]  <= 32'b	00011001110011101100100101111000	;
		random_num_table[148]  <= 32'b	00001111100101010101010100110011	;
		random_num_table[149]  <= 32'b	00010110011000010111000001011101	;
		random_num_table[150]  <= 32'b	00011000111011100000001001001110	;
		random_num_table[151]  <= 32'b	00001100001011001000011011011100	;
		random_num_table[152]  <= 32'b	00000011110000001011100011100111	;
		random_num_table[153]  <= 32'b	00000001011001100110111000001101	;
		random_num_table[154]  <= 32'b	00000100001000101101000001110101	;
		random_num_table[155]  <= 32'b	00010011000000101011010110000100	;
		random_num_table[156]  <= 32'b	00000100000011011000111100000111	;
		random_num_table[157]  <= 32'b	00011001010110010101110101100100	;
		random_num_table[158]  <= 32'b	00000101000101100111011101010100	;
		random_num_table[159]  <= 32'b	00001101010111101111110011111001	;
		random_num_table[160]  <= 32'b	00010101111010001001101000101110	;
		random_num_table[161]  <= 32'b	00001100011000110101011000111001	;
		random_num_table[162]  <= 32'b	00011100011101010111100100111111	;
		random_num_table[163]  <= 32'b	00011010110111000111000101000110	;
		random_num_table[164]  <= 32'b	00001101100111010000010100010011	;
		random_num_table[165]  <= 32'b	00010100010101011100000010000111	;
		random_num_table[166]  <= 32'b	00001010100010000101111100111100	;
		random_num_table[167]  <= 32'b	00000000110111000111010111110111	;
		random_num_table[168]  <= 32'b	00010111000100100011101101001100	;
		random_num_table[169]  <= 32'b	00001000011100101100111011110110	;
		random_num_table[170]  <= 32'b	00001111010110111011001111010110	;
		random_num_table[171]  <= 32'b	00010000010011101010100111100001	;
		random_num_table[172]  <= 32'b	00011011000110101000011010100010	;
		random_num_table[173]  <= 32'b	00001110100010110000100011111100	;
		random_num_table[174]  <= 32'b	00010101110000010111010010000100	;
		random_num_table[175]  <= 32'b	00010100011011111011110110101101	;
		random_num_table[176]  <= 32'b	00001110010101100100101101100111	;
		random_num_table[177]  <= 32'b	00000111111101110101001101000001	;
		random_num_table[178]  <= 32'b	00011010010110101101100101010111	;
		random_num_table[179]  <= 32'b	00000001111000011011001000110011	;
		random_num_table[180]  <= 32'b	00001100001000111011111001101000	;
		random_num_table[181]  <= 32'b	00010000100100101011100001110010	;
		random_num_table[182]  <= 32'b	00011000101111011011010100101100	;
		random_num_table[183]  <= 32'b	00001011000000110110110001001001	;
		random_num_table[184]  <= 32'b	00010110101001101111111101111000	;
		random_num_table[185]  <= 32'b	00010101011001101100100000110111	;
		random_num_table[186]  <= 32'b	00011100111000100010111010110011	;
		random_num_table[187]  <= 32'b	00011100010000101010110110010101	;
		random_num_table[188]  <= 32'b	00001110111110000111101111001011	;
		random_num_table[189]  <= 32'b	00010101100111010011111011000001	;
		random_num_table[190]  <= 32'b	00011011010110111010010101000111	;
		random_num_table[191]  <= 32'b	00010010100001110110100011111010	;
		random_num_table[192]  <= 32'b	00001001100110101101111010000001	;
		random_num_table[193]  <= 32'b	00011010110101001001010011100010	;
		random_num_table[194]  <= 32'b	00011000000011001111111110010011	;
		random_num_table[195]  <= 32'b	00010111101100010111010001010011	;
		random_num_table[196]  <= 32'b	00000111001100101100100101011101	;
		random_num_table[197]  <= 32'b	00000111011111011100111000110110	;
		random_num_table[198]  <= 32'b	00000000111111100011100110110110	;
		random_num_table[199]  <= 32'b	00010000000001000001010110100001	;
		random_num_table[200]  <= 32'b	00010101011011110111011110101000	;
		random_num_table[201]  <= 32'b	00001001100101100101000001011110	;
		random_num_table[202]  <= 32'b	00000010000001101001110011100111	;
		random_num_table[203]  <= 32'b	00010011111011100011111011011101	;
		random_num_table[204]  <= 32'b	00000011011000100101001000001001	;
		random_num_table[205]  <= 32'b	00000101101100011110000001100011	;
		random_num_table[206]  <= 32'b	00011000000010101110110010001101	;
		random_num_table[207]  <= 32'b	00000010111111000011011000110111	;
		random_num_table[208]  <= 32'b	00000000111000111110001011011111	;
		random_num_table[209]  <= 32'b	00001010100010101110101111010110	;
		random_num_table[210]  <= 32'b	00001111101101101001001100011110	;
		random_num_table[211]  <= 32'b	00001101101010111110010001100100	;
		random_num_table[212]  <= 32'b	00001001001111101011100100011100	;
		random_num_table[213]  <= 32'b	00001000010010000110010000101101	;
		random_num_table[214]  <= 32'b	00001010010100000011110010101110	;
		random_num_table[215]  <= 32'b	00000101000101110000101100100111	;
		random_num_table[216]  <= 32'b	00011001111011001101100011111001	;
		random_num_table[217]  <= 32'b	00011110101010110000110000001111	;
		random_num_table[218]  <= 32'b	00000010010000100110011010100011	;
		random_num_table[219]  <= 32'b	00001011011101010010011101010001	;
		random_num_table[220]  <= 32'b	00001011101110001011111011001011	;
		random_num_table[221]  <= 32'b	00011110000100111101101111111001	;
		random_num_table[222]  <= 32'b	00010101100101100010001000100100	;
		random_num_table[223]  <= 32'b	00010111011010000110001011001001	;
		random_num_table[224]  <= 32'b	00010000100101110110111110100010	;
		random_num_table[225]  <= 32'b	00000001111100010011000001001101	;
		random_num_table[226]  <= 32'b	00011111010001100101100100111001	;
		random_num_table[227]  <= 32'b	00000100001110110101011100000010	;
		random_num_table[228]  <= 32'b	00010110000111001110101011011010	;
		random_num_table[229]  <= 32'b	00000111110101101111111001110010	;
		random_num_table[230]  <= 32'b	00011010100010110101000100010101	;
		random_num_table[231]  <= 32'b	00000001010011101111110111111000	;
		random_num_table[232]  <= 32'b	00000011100001001011011100111100	;
		random_num_table[233]  <= 32'b	00010010101000100000101110110000	;
		random_num_table[234]  <= 32'b	00001000010010011011010110110110	;
		random_num_table[235]  <= 32'b	00001001001010010111110101110101	;
		random_num_table[236]  <= 32'b	00001100001001011011000011001110	;
		random_num_table[237]  <= 32'b	00001100100001010101111010000000	;
		random_num_table[238]  <= 32'b	00011100110111011010011001000001	;
		random_num_table[239]  <= 32'b	00000010100000010110011010111010	;
		random_num_table[240]  <= 32'b	00001001001011100100000111111100	;
		random_num_table[241]  <= 32'b	00001010011100011110101001001111	;
		random_num_table[242]  <= 32'b	00010000001011011110110110000110	;
		random_num_table[243]  <= 32'b	00001111101100010101011101100010	;
		random_num_table[244]  <= 32'b	00001100011000110110100110010001	;
		random_num_table[245]  <= 32'b	00000110111000000010111101010000	;
		random_num_table[246]  <= 32'b	00011101101000010111000010000101	;
		random_num_table[247]  <= 32'b	00001001010001111010011011100111	;
		random_num_table[248]  <= 32'b	00010000110001010101101111011001	;
		random_num_table[249]  <= 32'b	00001100111110111010001110110000	;
		random_num_table[250]  <= 32'b	00011010001011100000100110111011	;
		random_num_table[251]  <= 32'b	00010111100111111101001011110000	;
		random_num_table[252]  <= 32'b	00011110110101010000101001111110	;
		random_num_table[253]  <= 32'b	00001000001001110101010101111000	;
		random_num_table[254]  <= 32'b	00010010010101110011011001101110	;
		random_num_table[255]  <= 32'b	00011110011100110100011011100001	;			
	end
endmodule
