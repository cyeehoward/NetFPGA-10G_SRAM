`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:54:50 01/19/2015 
// Design Name: 
// Module Name:    rand_table_7 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module rand_table_11(axi_aclk , axi_aresetn , index_num , rand_out , en);
	input			axi_aclk , axi_aresetn , en;
	input		[7:0]	index_num;
	output		[31:0]	rand_out;

	reg 		[31:0]	random_num_table  [255:0];

	assign rand_out = en?random_num_table[index_num]:32'd0;
	
	always@(posedge axi_aclk)
	begin
		random_num_table[0]  <= 32'b	00001000110001000111010111111000	;
		random_num_table[1]  <= 32'b	00010000000100101010000101100001	;
		random_num_table[2]  <= 32'b	00000101111000000100101000000010	;
		random_num_table[3]  <= 32'b	00011110010001110110000110011100	;
		random_num_table[4]  <= 32'b	00000010000101110001110000110110	;
		random_num_table[5]  <= 32'b	00000100001101010011111001001101	;
		random_num_table[6]  <= 32'b	00001101001100110000101101100001	;
		random_num_table[7]  <= 32'b	00000110010011000000001101000010	;
		random_num_table[8]  <= 32'b	00001100100100010101101011001001	;
		random_num_table[9]  <= 32'b	00000100011100100001000101110011	;
		random_num_table[10]  <= 32'b	00010000100010011000001110110101	;
		random_num_table[11]  <= 32'b	00000111001100110100010010110110	;
		random_num_table[12]  <= 32'b	00000100010100001011110110010100	;
		random_num_table[13]  <= 32'b	00011001011111000011101011011011	;
		random_num_table[14]  <= 32'b	00010101111001111110001010011001	;
		random_num_table[15]  <= 32'b	00011110111010101100000111001100	;
		random_num_table[16]  <= 32'b	00000000100100000100011110011000	;
		random_num_table[17]  <= 32'b	00011110011110111000000011001001	;
		random_num_table[18]  <= 32'b	00001101101000000110111101001111	;
		random_num_table[19]  <= 32'b	00010110111101101011110110001100	;
		random_num_table[20]  <= 32'b	00000000010000110101101111110100	;
		random_num_table[21]  <= 32'b	00001011101011101110110101011001	;
		random_num_table[22]  <= 32'b	00001101001011100001000011111111	;
		random_num_table[23]  <= 32'b	00000011110100111101010110011110	;
		random_num_table[24]  <= 32'b	00000101101011110111001101110011	;
		random_num_table[25]  <= 32'b	00010010000101010101111010100010	;
		random_num_table[26]  <= 32'b	00010100101100100111011111110011	;
		random_num_table[27]  <= 32'b	00001010001111011011110100000100	;
		random_num_table[28]  <= 32'b	00010010000111010000011010101110	;
		random_num_table[29]  <= 32'b	00000111010101111110110001111001	;
		random_num_table[30]  <= 32'b	00001110010110100010110101001000	;
		random_num_table[31]  <= 32'b	00011001101111100110000010011110	;
		random_num_table[32]  <= 32'b	00010001101101001110100000110101	;
		random_num_table[33]  <= 32'b	00001111001100010010101000100110	;
		random_num_table[34]  <= 32'b	00011100011001000011011111000101	;
		random_num_table[35]  <= 32'b	00010101110001100001000101010100	;
		random_num_table[36]  <= 32'b	00000001111100000011011100000111	;
		random_num_table[37]  <= 32'b	00001010010101100011110111100110	;
		random_num_table[38]  <= 32'b	00010101000001010010001010111010	;
		random_num_table[39]  <= 32'b	00001111101010101111000101111111	;
		random_num_table[40]  <= 32'b	00000101000111000001110011010111	;
		random_num_table[41]  <= 32'b	00011010101011000101111110110100	;
		random_num_table[42]  <= 32'b	00000001010000011101111000101101	;
		random_num_table[43]  <= 32'b	00001010001010010011111000111001	;
		random_num_table[44]  <= 32'b	00011011110011011111111001010110	;
		random_num_table[45]  <= 32'b	00000001101000101011000001101101	;
		random_num_table[46]  <= 32'b	00000110000100000010000011110001	;
		random_num_table[47]  <= 32'b	00001011100011110110010001011000	;
		random_num_table[48]  <= 32'b	00011101100001001100110010110110	;
		random_num_table[49]  <= 32'b	00000111101110110111011110000001	;
		random_num_table[50]  <= 32'b	00001100001100000100100101001111	;
		random_num_table[51]  <= 32'b	00000001010011001101100000010110	;
		random_num_table[52]  <= 32'b	00000000001001100110010011001001	;
		random_num_table[53]  <= 32'b	00001010001011000001001010100001	;
		random_num_table[54]  <= 32'b	00011001011100100110111001001001	;
		random_num_table[55]  <= 32'b	00000001101101011110011011001010	;
		random_num_table[56]  <= 32'b	00011100100001110010001001110010	;
		random_num_table[57]  <= 32'b	00001000100000001011100111011000	;
		random_num_table[58]  <= 32'b	00010110111111011111111001001110	;
		random_num_table[59]  <= 32'b	00001010011110110110110100100011	;
		random_num_table[60]  <= 32'b	00010001001110110001001100011010	;
		random_num_table[61]  <= 32'b	00000111000111001001010101010110	;
		random_num_table[62]  <= 32'b	00011110110110100100101011010010	;
		random_num_table[63]  <= 32'b	00001000111100110100010100001010	;
		random_num_table[64]  <= 32'b	00011110000000101101000110100111	;
		random_num_table[65]  <= 32'b	00000000000000100010100111100011	;
		random_num_table[66]  <= 32'b	00010110111111001100110000111101	;
		random_num_table[67]  <= 32'b	00001011011001100011001001111001	;
		random_num_table[68]  <= 32'b	00010101111011011111000100010101	;
		random_num_table[69]  <= 32'b	00011011111011111100011100100101	;
		random_num_table[70]  <= 32'b	00001010011000011100110011101000	;
		random_num_table[71]  <= 32'b	00000110101011001110101101001001	;
		random_num_table[72]  <= 32'b	00001110010111110011110001111010	;
		random_num_table[73]  <= 32'b	00011001000001110110100010111011	;
		random_num_table[74]  <= 32'b	00010101001001010100011001110110	;
		random_num_table[75]  <= 32'b	00001010101001101011100100111011	;
		random_num_table[76]  <= 32'b	00000101010000010011101000101010	;
		random_num_table[77]  <= 32'b	00011111111001101101000110000000	;
		random_num_table[78]  <= 32'b	00010110000000101110000001101001	;
		random_num_table[79]  <= 32'b	00000101100001001001101010000101	;
		random_num_table[80]  <= 32'b	00001110001011100001100000100010	;
		random_num_table[81]  <= 32'b	00010010000100001101000011001111	;
		random_num_table[82]  <= 32'b	00011011101111100010001010101110	;
		random_num_table[83]  <= 32'b	00010000111101010110110111001100	;
		random_num_table[84]  <= 32'b	00001010011000110111111000010011	;
		random_num_table[85]  <= 32'b	00000011101101110000101101000010	;
		random_num_table[86]  <= 32'b	00000110001100111010001110010101	;
		random_num_table[87]  <= 32'b	00001011110111111110110111010100	;
		random_num_table[88]  <= 32'b	00011101101011101100011110101011	;
		random_num_table[89]  <= 32'b	00000011111011010101100110011011	;
		random_num_table[90]  <= 32'b	00010110000010001000010011100110	;
		random_num_table[91]  <= 32'b	00011111111000101100101110011010	;
		random_num_table[92]  <= 32'b	00011001111100100100110111100101	;
		random_num_table[93]  <= 32'b	00011100111001000011101111011000	;
		random_num_table[94]  <= 32'b	00000000111111000100111000010001	;
		random_num_table[95]  <= 32'b	00010010001011110101100100100001	;
		random_num_table[96]  <= 32'b	00011010111100001110101001100111	;
		random_num_table[97]  <= 32'b	00011000100000101010010011111000	;
		random_num_table[98]  <= 32'b	00010100100110011100011101100010	;
		random_num_table[99]  <= 32'b	00011101010011111010001100001101	;
		random_num_table[100]  <= 32'b	00001010010011011110001110111110	;
		random_num_table[101]  <= 32'b	00010101001000100100011101011110	;
		random_num_table[102]  <= 32'b	00010101010010111010010010111111	;
		random_num_table[103]  <= 32'b	00001010110101000101100111110110	;
		random_num_table[104]  <= 32'b	00010111000100010011011011001000	;
		random_num_table[105]  <= 32'b	00001101000111000111101011011000	;
		random_num_table[106]  <= 32'b	00010011010111011000101010000000	;
		random_num_table[107]  <= 32'b	00000001110010110001001010011111	;
		random_num_table[108]  <= 32'b	00000101101110100010101000011110	;
		random_num_table[109]  <= 32'b	00010111101000110010100000000111	;
		random_num_table[110]  <= 32'b	00001011110111101100111111101101	;
		random_num_table[111]  <= 32'b	00010110011100000010010110010101	;
		random_num_table[112]  <= 32'b	00011100001011011110100110010110	;
		random_num_table[113]  <= 32'b	00010001001111100101001010000100	;
		random_num_table[114]  <= 32'b	00001110110101100011001110111101	;
		random_num_table[115]  <= 32'b	00010100010001010000010110110011	;
		random_num_table[116]  <= 32'b	00010000000111000111110111111010	;
		random_num_table[117]  <= 32'b	00010011110100111100101111001101	;
		random_num_table[118]  <= 32'b	00001111100111100101010110110110	;
		random_num_table[119]  <= 32'b	00001010001001111110010110010000	;
		random_num_table[120]  <= 32'b	00010001101111111111011110110001	;
		random_num_table[121]  <= 32'b	00011101110011011100110010111110	;
		random_num_table[122]  <= 32'b	00010010011010010100000101000010	;
		random_num_table[123]  <= 32'b	00011010010001100111010000001000	;
		random_num_table[124]  <= 32'b	00011101010010001000011000000001	;
		random_num_table[125]  <= 32'b	00001001011100110111111001010001	;
		random_num_table[126]  <= 32'b	00000011010011000000011001110101	;
		random_num_table[127]  <= 32'b	00000111100111001110100111101111	;
		random_num_table[128]  <= 32'b	00001001101100110011101011100000	;
		random_num_table[129]  <= 32'b	00011101011001110010000101101001	;
		random_num_table[130]  <= 32'b	00000111001010100111101110101000	;
		random_num_table[131]  <= 32'b	00001000010000101110111110001101	;
		random_num_table[132]  <= 32'b	00000110010110010100011101110001	;
		random_num_table[133]  <= 32'b	00010100000011000111101110011011	;
		random_num_table[134]  <= 32'b	00000001011101011001001111111010	;
		random_num_table[135]  <= 32'b	00010111000001010000111110011100	;
		random_num_table[136]  <= 32'b	00001111001010010100000001001110	;
		random_num_table[137]  <= 32'b	00010111001110110111010001000001	;
		random_num_table[138]  <= 32'b	00001110011011001101001001000101	;
		random_num_table[139]  <= 32'b	00011101110000001101101000010000	;
		random_num_table[140]  <= 32'b	00000000101101111110000101100110	;
		random_num_table[141]  <= 32'b	00011111101111000110010001001111	;
		random_num_table[142]  <= 32'b	00011101101111000101001000011011	;
		random_num_table[143]  <= 32'b	00001011110010111010010000101011	;
		random_num_table[144]  <= 32'b	00010011101101111110101111110001	;
		random_num_table[145]  <= 32'b	00010110101011000000000101000010	;
		random_num_table[146]  <= 32'b	00000010000010010001011100110000	;
		random_num_table[147]  <= 32'b	00011101100010001000101110110001	;
		random_num_table[148]  <= 32'b	00011000101011101001110011010101	;
		random_num_table[149]  <= 32'b	00010010100101101001010010000001	;
		random_num_table[150]  <= 32'b	00011101100111001010011000100101	;
		random_num_table[151]  <= 32'b	00001011110110101001100011110110	;
		random_num_table[152]  <= 32'b	00000110111010110010110011111100	;
		random_num_table[153]  <= 32'b	00000011111101010010101001111111	;
		random_num_table[154]  <= 32'b	00001111011101001111101111110001	;
		random_num_table[155]  <= 32'b	00001001101111110001110110001110	;
		random_num_table[156]  <= 32'b	00011000010011100011110111100110	;
		random_num_table[157]  <= 32'b	00010011010111001111101011001001	;
		random_num_table[158]  <= 32'b	00010010111101000101110111101110	;
		random_num_table[159]  <= 32'b	00000001011101111111100000000000	;
		random_num_table[160]  <= 32'b	00001001000101111100101110101111	;
		random_num_table[161]  <= 32'b	00011101010111011011101100101010	;
		random_num_table[162]  <= 32'b	00001001100010011110101001000001	;
		random_num_table[163]  <= 32'b	00000000111101100011000011001111	;
		random_num_table[164]  <= 32'b	00010111100010011000011100110100	;
		random_num_table[165]  <= 32'b	00010110111100111110110101100110	;
		random_num_table[166]  <= 32'b	00000001000101001001011011110001	;
		random_num_table[167]  <= 32'b	00011011011000100001101100111010	;
		random_num_table[168]  <= 32'b	00001001001101011100001101111110	;
		random_num_table[169]  <= 32'b	00010100101010001010001110000110	;
		random_num_table[170]  <= 32'b	00000111111010111010110001010100	;
		random_num_table[171]  <= 32'b	00011011001111110011000001100011	;
		random_num_table[172]  <= 32'b	00000011111010101111001011111000	;
		random_num_table[173]  <= 32'b	00000110011101110000100010110010	;
		random_num_table[174]  <= 32'b	00001010100110100110011110010011	;
		random_num_table[175]  <= 32'b	00001001001101011010101100111101	;
		random_num_table[176]  <= 32'b	00010110001000100110101010010011	;
		random_num_table[177]  <= 32'b	00010111011010011101111110111011	;
		random_num_table[178]  <= 32'b	00011000110000000110001100010000	;
		random_num_table[179]  <= 32'b	00011010111110100011000000101100	;
		random_num_table[180]  <= 32'b	00001000110011010011000010011000	;
		random_num_table[181]  <= 32'b	00010001001001100011001011000011	;
		random_num_table[182]  <= 32'b	00001011111011100100110101111000	;
		random_num_table[183]  <= 32'b	00010000010101010010011111111000	;
		random_num_table[184]  <= 32'b	00010111011101011000011000111110	;
		random_num_table[185]  <= 32'b	00000111010101000010011001110000	;
		random_num_table[186]  <= 32'b	00010111011000001001001001101110	;
		random_num_table[187]  <= 32'b	00000011011000101111110101001111	;
		random_num_table[188]  <= 32'b	00011000110001110001010100100101	;
		random_num_table[189]  <= 32'b	00000111001100110010100101110010	;
		random_num_table[190]  <= 32'b	00011110011001110011011010010111	;
		random_num_table[191]  <= 32'b	00000111100101011101000011100111	;
		random_num_table[192]  <= 32'b	00011001101001000110100110111110	;
		random_num_table[193]  <= 32'b	00001000001011001010000101101110	;
		random_num_table[194]  <= 32'b	00011111010111010000111011001010	;
		random_num_table[195]  <= 32'b	00011000011110000011010010001001	;
		random_num_table[196]  <= 32'b	00001101100110000010010110010100	;
		random_num_table[197]  <= 32'b	00011000101011110011100010110011	;
		random_num_table[198]  <= 32'b	00000101000101100101010111111010	;
		random_num_table[199]  <= 32'b	00000000000110010101111001101010	;
		random_num_table[200]  <= 32'b	00011100111110011111000001100010	;
		random_num_table[201]  <= 32'b	00011000111010000111011111111010	;
		random_num_table[202]  <= 32'b	00011110110010101000011100100001	;
		random_num_table[203]  <= 32'b	00001001111111101111000010010100	;
		random_num_table[204]  <= 32'b	00001101110111110000000111101000	;
		random_num_table[205]  <= 32'b	00000101101001100101101011010010	;
		random_num_table[206]  <= 32'b	00010010011001100101001001110010	;
		random_num_table[207]  <= 32'b	00011111111100110111010110011001	;
		random_num_table[208]  <= 32'b	00010001111010010000100010101110	;
		random_num_table[209]  <= 32'b	00011110000111101011110111010001	;
		random_num_table[210]  <= 32'b	00010001110110010010111011000111	;
		random_num_table[211]  <= 32'b	00011111011100011110100000000011	;
		random_num_table[212]  <= 32'b	00000001111000010100111111111110	;
		random_num_table[213]  <= 32'b	00011100101100010011110110110011	;
		random_num_table[214]  <= 32'b	00000101010110111010100101111100	;
		random_num_table[215]  <= 32'b	00000101010101011000000100111101	;
		random_num_table[216]  <= 32'b	00001110101100001110010101001111	;
		random_num_table[217]  <= 32'b	00011110110110011001000011011100	;
		random_num_table[218]  <= 32'b	00010101011100001101110101011000	;
		random_num_table[219]  <= 32'b	00001100010110110101111011010111	;
		random_num_table[220]  <= 32'b	00000100101010001110101100100010	;
		random_num_table[221]  <= 32'b	00001001101011000110110100111001	;
		random_num_table[222]  <= 32'b	00000100101011000001000101111101	;
		random_num_table[223]  <= 32'b	00000011111010101110000101001101	;
		random_num_table[224]  <= 32'b	00011000011111001110111111101111	;
		random_num_table[225]  <= 32'b	00000011010011000110011000111101	;
		random_num_table[226]  <= 32'b	00010100100111111100000111110001	;
		random_num_table[227]  <= 32'b	00011100110111100000101110100001	;
		random_num_table[228]  <= 32'b	00000111010000001111111110110101	;
		random_num_table[229]  <= 32'b	00001100011110110110101110101101	;
		random_num_table[230]  <= 32'b	00001001011001100111100001101101	;
		random_num_table[231]  <= 32'b	00010110010001100110001011010000	;
		random_num_table[232]  <= 32'b	00000011011100001001000101101010	;
		random_num_table[233]  <= 32'b	00010101111100010111111111011010	;
		random_num_table[234]  <= 32'b	00011111101010111001010100000010	;
		random_num_table[235]  <= 32'b	00000110000010100111101011000101	;
		random_num_table[236]  <= 32'b	00000100010011000010100110111001	;
		random_num_table[237]  <= 32'b	00011011000100010011011101001101	;
		random_num_table[238]  <= 32'b	00001010011100101100000010101101	;
		random_num_table[239]  <= 32'b	00001011000000101100101101111111	;
		random_num_table[240]  <= 32'b	00010001001010010101011011100101	;
		random_num_table[241]  <= 32'b	00010010110101010000111100010101	;
		random_num_table[242]  <= 32'b	00000001001000110110001110000000	;
		random_num_table[243]  <= 32'b	00010111010010101100011010111011	;
		random_num_table[244]  <= 32'b	00000100100001011010101000100110	;
		random_num_table[245]  <= 32'b	00010110001011001011100110001110	;
		random_num_table[246]  <= 32'b	00000111000001010110011100001110	;
		random_num_table[247]  <= 32'b	00001111001001000100010100101111	;
		random_num_table[248]  <= 32'b	00011001001000000110000110100110	;
		random_num_table[249]  <= 32'b	00011101111010100010111011001101	;
		random_num_table[250]  <= 32'b	00001101000111100110111000000100	;
		random_num_table[251]  <= 32'b	00001011000100110101010010111100	;
		random_num_table[252]  <= 32'b	00011110100010100011001110101101	;
		random_num_table[253]  <= 32'b	00011011100010111101100010111101	;
		random_num_table[254]  <= 32'b	00010010100010000111101110100100	;
		random_num_table[255]  <= 32'b	00001110110101101010111010000001	;			
	end
endmodule
