`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:51:43 01/19/2015 
// Design Name: 
// Module Name:    rand_table_2 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module rand_table_2(axi_aclk , axi_aresetn , index_num , rand_out , en);
	input			axi_aclk , axi_aresetn , en;
	input		[7:0]	index_num;
	output		[31:0]	rand_out;

	reg 		[31:0]	random_num_table  [255:0];

	assign rand_out = en?random_num_table[index_num]:32'd0;
	
	always@(posedge axi_aclk)
	begin
		random_num_table[0]  <= 32'b	00011010011111100001000001011011	;
		random_num_table[1]  <= 32'b	00011010011010001000101011110001	;
		random_num_table[2]  <= 32'b	00001110001001110110101000111011	;
		random_num_table[3]  <= 32'b	00010110110000001001111010001110	;
		random_num_table[4]  <= 32'b	00000001010101011110001000011000	;
		random_num_table[5]  <= 32'b	00001110010000011100010010101000	;
		random_num_table[6]  <= 32'b	00001101101110100000110110010101	;
		random_num_table[7]  <= 32'b	00010001100110010110001101001101	;
		random_num_table[8]  <= 32'b	00000000000100111111000110011001	;
		random_num_table[9]  <= 32'b	00010110110111010101001011001101	;
		random_num_table[10]  <= 32'b	00001011100111011001101010110100	;
		random_num_table[11]  <= 32'b	00010111001010001010101110011101	;
		random_num_table[12]  <= 32'b	00011100110101001110000100100100	;
		random_num_table[13]  <= 32'b	00011001101011111111110011101011	;
		random_num_table[14]  <= 32'b	00010001011110111110001010111010	;
		random_num_table[15]  <= 32'b	00001100111100010010001010010111	;
		random_num_table[16]  <= 32'b	00000010111111010110101000111110	;
		random_num_table[17]  <= 32'b	00001101111101001001011000010001	;
		random_num_table[18]  <= 32'b	00000000011110100110011001101110	;
		random_num_table[19]  <= 32'b	00000101010101011010010101101000	;
		random_num_table[20]  <= 32'b	00010101010011101110011100001001	;
		random_num_table[21]  <= 32'b	00010011000001001000110000100111	;
		random_num_table[22]  <= 32'b	00001110101111011110011000101011	;
		random_num_table[23]  <= 32'b	00000101100100001100101101111011	;
		random_num_table[24]  <= 32'b	00011000100001010111101000111000	;
		random_num_table[25]  <= 32'b	00011000010000101011010111010101	;
		random_num_table[26]  <= 32'b	00010101101110010100011101000101	;
		random_num_table[27]  <= 32'b	00011111100010101000001110010100	;
		random_num_table[28]  <= 32'b	00000001001001110100010100100110	;
		random_num_table[29]  <= 32'b	00000000011000011101010011101000	;
		random_num_table[30]  <= 32'b	00010101101101010010001111110010	;
		random_num_table[31]  <= 32'b	00011000101110011010010000010101	;
		random_num_table[32]  <= 32'b	00011110110100011111111110110101	;
		random_num_table[33]  <= 32'b	00000001011101100100101100010011	;
		random_num_table[34]  <= 32'b	00011101010100011111001101111101	;
		random_num_table[35]  <= 32'b	00011110000110100110101001101000	;
		random_num_table[36]  <= 32'b	00010011010011000001100010111001	;
		random_num_table[37]  <= 32'b	00001001011110101011000111010011	;
		random_num_table[38]  <= 32'b	00010101100010000100101100111110	;
		random_num_table[39]  <= 32'b	00010000010001101100011101010111	;
		random_num_table[40]  <= 32'b	00010000101111001110001011001110	;
		random_num_table[41]  <= 32'b	00001011110000100001110011110110	;
		random_num_table[42]  <= 32'b	00001101011100100111000100011111	;
		random_num_table[43]  <= 32'b	00001001010000001010101111000010	;
		random_num_table[44]  <= 32'b	00000110001010000000100101011110	;
		random_num_table[45]  <= 32'b	00001010010111110000101111011001	;
		random_num_table[46]  <= 32'b	00001101010000000000010001001011	;
		random_num_table[47]  <= 32'b	00001000011101111100100001100100	;
		random_num_table[48]  <= 32'b	00001100000011011111001110111101	;
		random_num_table[49]  <= 32'b	00010011101101110000111000011111	;
		random_num_table[50]  <= 32'b	00001100001001010010101000101011	;
		random_num_table[51]  <= 32'b	00010111001110111111001101000001	;
		random_num_table[52]  <= 32'b	00001000011010001100001011010000	;
		random_num_table[53]  <= 32'b	00010000011010011111101100001110	;
		random_num_table[54]  <= 32'b	00011010001110111011101110010111	;
		random_num_table[55]  <= 32'b	00011110101100010001110011100011	;
		random_num_table[56]  <= 32'b	00010101111001101011101111000101	;
		random_num_table[57]  <= 32'b	00001001001111110101100110011111	;
		random_num_table[58]  <= 32'b	00010011110100111011100001010110	;
		random_num_table[59]  <= 32'b	00010001100110001000011010001111	;
		random_num_table[60]  <= 32'b	00010010100000011110001101011100	;
		random_num_table[61]  <= 32'b	00000111100000000001010011010111	;
		random_num_table[62]  <= 32'b	00000011100001100111111011011111	;
		random_num_table[63]  <= 32'b	00000011111000000010011001111010	;
		random_num_table[64]  <= 32'b	00000001011010001111011011111110	;
		random_num_table[65]  <= 32'b	00000010000110000110010011000100	;
		random_num_table[66]  <= 32'b	00011111110101001101110000000001	;
		random_num_table[67]  <= 32'b	00001111101101011011100111011000	;
		random_num_table[68]  <= 32'b	00011101010100001111001011000000	;
		random_num_table[69]  <= 32'b	00001011010111111000111110011101	;
		random_num_table[70]  <= 32'b	00011100101010001010100011100001	;
		random_num_table[71]  <= 32'b	00010011111011001110010011010111	;
		random_num_table[72]  <= 32'b	00000111110111100001110010010001	;
		random_num_table[73]  <= 32'b	00010001111000110110101001111000	;
		random_num_table[74]  <= 32'b	00000001010101100011100010011000	;
		random_num_table[75]  <= 32'b	00011110100100000100101011110000	;
		random_num_table[76]  <= 32'b	00011111010000110111111011111101	;
		random_num_table[77]  <= 32'b	00001001001101101011010001010101	;
		random_num_table[78]  <= 32'b	00000010100011100100011110011100	;
		random_num_table[79]  <= 32'b	00010010111001110101100111010000	;
		random_num_table[80]  <= 32'b	00010010001001010010100100010100	;
		random_num_table[81]  <= 32'b	00000001101000101111000100110000	;
		random_num_table[82]  <= 32'b	00001111010111100011001001111000	;
		random_num_table[83]  <= 32'b	00010010000111011001110010001011	;
		random_num_table[84]  <= 32'b	00001111001010101011110010111001	;
		random_num_table[85]  <= 32'b	00010110001010101011101101100110	;
		random_num_table[86]  <= 32'b	00000110010101011010100111010110	;
		random_num_table[87]  <= 32'b	00011111000101100110110101001111	;
		random_num_table[88]  <= 32'b	00010011100111010010000111000010	;
		random_num_table[89]  <= 32'b	00010000001010011100101111010010	;
		random_num_table[90]  <= 32'b	00001111010011110100100011111100	;
		random_num_table[91]  <= 32'b	00000010011011000100100101000010	;
		random_num_table[92]  <= 32'b	00000100011011001001110001101101	;
		random_num_table[93]  <= 32'b	00010111111010000100110010001011	;
		random_num_table[94]  <= 32'b	00001111010010100001110001110110	;
		random_num_table[95]  <= 32'b	00010001011000000010000111111101	;
		random_num_table[96]  <= 32'b	00001101000111000000010100011110	;
		random_num_table[97]  <= 32'b	00000100100100110110010010100111	;
		random_num_table[98]  <= 32'b	00000001111000101110100011001111	;
		random_num_table[99]  <= 32'b	00000101110111111101101010000111	;
		random_num_table[100]  <= 32'b	00000000101101011100110110111000	;
		random_num_table[101]  <= 32'b	00011000011011101111010111010001	;
		random_num_table[102]  <= 32'b	00011110011101111001011100100110	;
		random_num_table[103]  <= 32'b	00001001001101111000011110101000	;
		random_num_table[104]  <= 32'b	00000110010100001001001111100011	;
		random_num_table[105]  <= 32'b	00011111000101100101000111100001	;
		random_num_table[106]  <= 32'b	00000110000101001001100111101001	;
		random_num_table[107]  <= 32'b	00011011001111111111000101000111	;
		random_num_table[108]  <= 32'b	00000100100101111111000100111000	;
		random_num_table[109]  <= 32'b	00010110111101000111110011010011	;
		random_num_table[110]  <= 32'b	00001111011011101000010110010100	;
		random_num_table[111]  <= 32'b	00010110100111100110000110010100	;
		random_num_table[112]  <= 32'b	00011110010001100111101010001100	;
		random_num_table[113]  <= 32'b	00001011010101010001101111010010	;
		random_num_table[114]  <= 32'b	00011011111110111001011111111111	;
		random_num_table[115]  <= 32'b	00001110001010001100111101010001	;
		random_num_table[116]  <= 32'b	00010011011011100001001010011110	;
		random_num_table[117]  <= 32'b	00010010011110001000001100011100	;
		random_num_table[118]  <= 32'b	00011000110010010100110110010000	;
		random_num_table[119]  <= 32'b	00010000111101111010010011011010	;
		random_num_table[120]  <= 32'b	00010100101000001100010001011011	;
		random_num_table[121]  <= 32'b	00000011010011101100111101011101	;
		random_num_table[122]  <= 32'b	00000101100111101011110011010000	;
		random_num_table[123]  <= 32'b	00000101001001010010011011011010	;
		random_num_table[124]  <= 32'b	00000010110010100100000110010100	;
		random_num_table[125]  <= 32'b	00001100111111100001000001001000	;
		random_num_table[126]  <= 32'b	00010001111000110101101010110011	;
		random_num_table[127]  <= 32'b	00001101110100011011010011001100	;
		random_num_table[128]  <= 32'b	00011010001000110100110010010000	;
		random_num_table[129]  <= 32'b	00011001010100001011101110011000	;
		random_num_table[130]  <= 32'b	00000000110111111101010011010001	;
		random_num_table[131]  <= 32'b	00010000000110100111001101110010	;
		random_num_table[132]  <= 32'b	00001000110101001100111001001010	;
		random_num_table[133]  <= 32'b	00010101010101101100100101100011	;
		random_num_table[134]  <= 32'b	00010001100001110010001011000000	;
		random_num_table[135]  <= 32'b	00000100101111011011101011011100	;
		random_num_table[136]  <= 32'b	00010000000011011010010011000100	;
		random_num_table[137]  <= 32'b	00010000001000010101100010100000	;
		random_num_table[138]  <= 32'b	00001110111001101001011010111101	;
		random_num_table[139]  <= 32'b	00001100001100011010101000110010	;
		random_num_table[140]  <= 32'b	00010111110010000001001101011011	;
		random_num_table[141]  <= 32'b	00000000001010011001110001011111	;
		random_num_table[142]  <= 32'b	00010000110100000110110010110100	;
		random_num_table[143]  <= 32'b	00001011000010000001110110101010	;
		random_num_table[144]  <= 32'b	00001111000101101111010010010010	;
		random_num_table[145]  <= 32'b	00010110001111111011111010100000	;
		random_num_table[146]  <= 32'b	00000011001101000011000010000001	;
		random_num_table[147]  <= 32'b	00010101101100011011000101001001	;
		random_num_table[148]  <= 32'b	00011011000110000100110100101010	;
		random_num_table[149]  <= 32'b	00000100110011101011110001101101	;
		random_num_table[150]  <= 32'b	00011000110001111110011101100011	;
		random_num_table[151]  <= 32'b	00010011000001101011100000011010	;
		random_num_table[152]  <= 32'b	00001000000110110100001000010111	;
		random_num_table[153]  <= 32'b	00000010110000011101111101101010	;
		random_num_table[154]  <= 32'b	00011100011010011110110010101011	;
		random_num_table[155]  <= 32'b	00010110001010110111111000000100	;
		random_num_table[156]  <= 32'b	00010001100010010010111010100101	;
		random_num_table[157]  <= 32'b	00001010100001111101011101110001	;
		random_num_table[158]  <= 32'b	00001011110110100010001100100110	;
		random_num_table[159]  <= 32'b	00000111111101111110100101000110	;
		random_num_table[160]  <= 32'b	00010000010111111110011011010010	;
		random_num_table[161]  <= 32'b	00001110101110001011000100110101	;
		random_num_table[162]  <= 32'b	00011000010111010100100110100101	;
		random_num_table[163]  <= 32'b	00011011111111010111111011001011	;
		random_num_table[164]  <= 32'b	00011011000100011100111001010001	;
		random_num_table[165]  <= 32'b	00010001001110111101000001101101	;
		random_num_table[166]  <= 32'b	00001101011010111101011101101011	;
		random_num_table[167]  <= 32'b	00000110000111111100110101100001	;
		random_num_table[168]  <= 32'b	00001101011000100101000010110010	;
		random_num_table[169]  <= 32'b	00001011110100010001101111101100	;
		random_num_table[170]  <= 32'b	00011001110101011001010111010010	;
		random_num_table[171]  <= 32'b	00000111001110000010011001001100	;
		random_num_table[172]  <= 32'b	00000100001010001010111111101010	;
		random_num_table[173]  <= 32'b	00010011010010101001111011010001	;
		random_num_table[174]  <= 32'b	00001010100111001010000111110110	;
		random_num_table[175]  <= 32'b	00001010010001111111011110010110	;
		random_num_table[176]  <= 32'b	00000011100010011000110010010001	;
		random_num_table[177]  <= 32'b	00001000111101010111111101110111	;
		random_num_table[178]  <= 32'b	00001101011101001111000110111011	;
		random_num_table[179]  <= 32'b	00010000101010010101101110101100	;
		random_num_table[180]  <= 32'b	00010000001100000000110111101001	;
		random_num_table[181]  <= 32'b	00000011001010100011100010001000	;
		random_num_table[182]  <= 32'b	00011010010000101000111010001010	;
		random_num_table[183]  <= 32'b	00010011001000100100001000111101	;
		random_num_table[184]  <= 32'b	00010011000010011011110101110000	;
		random_num_table[185]  <= 32'b	00010101000010001000101100001110	;
		random_num_table[186]  <= 32'b	00011111110001000001001001111001	;
		random_num_table[187]  <= 32'b	00011010101110100010010011101110	;
		random_num_table[188]  <= 32'b	00001010000111010010101110111100	;
		random_num_table[189]  <= 32'b	00011111001110100010100001111010	;
		random_num_table[190]  <= 32'b	00001110111110001000000011001111	;
		random_num_table[191]  <= 32'b	00000101010001111000110010101111	;
		random_num_table[192]  <= 32'b	00010111011010101101011010000010	;
		random_num_table[193]  <= 32'b	00011111000010101111100010010110	;
		random_num_table[194]  <= 32'b	00010111100101111100001001100100	;
		random_num_table[195]  <= 32'b	00001000010010110010111001110000	;
		random_num_table[196]  <= 32'b	00000001001001100101000000101101	;
		random_num_table[197]  <= 32'b	00000100001110010101110011011100	;
		random_num_table[198]  <= 32'b	00010001001000111111010010001100	;
		random_num_table[199]  <= 32'b	00001111111101101111011101101110	;
		random_num_table[200]  <= 32'b	00010000111110010100100110111100	;
		random_num_table[201]  <= 32'b	00010001001100110011101111011001	;
		random_num_table[202]  <= 32'b	00010000011010101100100010100101	;
		random_num_table[203]  <= 32'b	00011010101101100000011001100000	;
		random_num_table[204]  <= 32'b	00001001011101100001101111101111	;
		random_num_table[205]  <= 32'b	00001101010000110111111111100000	;
		random_num_table[206]  <= 32'b	00010001001100000001000100110010	;
		random_num_table[207]  <= 32'b	00010110110100101001100100101111	;
		random_num_table[208]  <= 32'b	00000100100001110000000000000010	;
		random_num_table[209]  <= 32'b	00001101001111101011010100100010	;
		random_num_table[210]  <= 32'b	00010010110011010001110100110101	;
		random_num_table[211]  <= 32'b	00011010100000100110100010000111	;
		random_num_table[212]  <= 32'b	00010110000111010101110001000110	;
		random_num_table[213]  <= 32'b	00011010100100110011101110101101	;
		random_num_table[214]  <= 32'b	00011100100000111110001100101011	;
		random_num_table[215]  <= 32'b	00001101010010001110010000101000	;
		random_num_table[216]  <= 32'b	00000010010101111001101010111110	;
		random_num_table[217]  <= 32'b	00010101011010001011110101101101	;
		random_num_table[218]  <= 32'b	00010100110100001100101111110011	;
		random_num_table[219]  <= 32'b	00000100100111000101000010111010	;
		random_num_table[220]  <= 32'b	00000000010111010100110011011101	;
		random_num_table[221]  <= 32'b	00001101001110011111000011101000	;
		random_num_table[222]  <= 32'b	00001110000110111110000101110001	;
		random_num_table[223]  <= 32'b	00000000111001011111011011011101	;
		random_num_table[224]  <= 32'b	00011111111011101100100111111000	;
		random_num_table[225]  <= 32'b	00011111010101011001101001001001	;
		random_num_table[226]  <= 32'b	00001000110001010000110010100011	;
		random_num_table[227]  <= 32'b	00010001111011010010010111100111	;
		random_num_table[228]  <= 32'b	00011011001111110101001100101111	;
		random_num_table[229]  <= 32'b	00010101001001000000001101101010	;
		random_num_table[230]  <= 32'b	00001000111011111110011001111011	;
		random_num_table[231]  <= 32'b	00011111111010110101110010010001	;
		random_num_table[232]  <= 32'b	00010011001001001010010101011010	;
		random_num_table[233]  <= 32'b	00011101011111011001100011011101	;
		random_num_table[234]  <= 32'b	00000111010011101111110010100110	;
		random_num_table[235]  <= 32'b	00010011111101101010101101110001	;
		random_num_table[236]  <= 32'b	00000001110100000000101110101000	;
		random_num_table[237]  <= 32'b	00001101001000100001101000001100	;
		random_num_table[238]  <= 32'b	00010000010011111111000101110000	;
		random_num_table[239]  <= 32'b	00000011000010111111100101101000	;
		random_num_table[240]  <= 32'b	00011011001101010001110010010010	;
		random_num_table[241]  <= 32'b	00001000100101000000011010011101	;
		random_num_table[242]  <= 32'b	00001111011001111000010001101011	;
		random_num_table[243]  <= 32'b	00010101110011001001111010101110	;
		random_num_table[244]  <= 32'b	00011101101110001011000001001100	;
		random_num_table[245]  <= 32'b	00011001001111001000111110101100	;
		random_num_table[246]  <= 32'b	00010001111001001100011001011111	;
		random_num_table[247]  <= 32'b	00010000011101010110000000101000	;
		random_num_table[248]  <= 32'b	00001101010101010100011010101101	;
		random_num_table[249]  <= 32'b	00001111100110100001110101001101	;
		random_num_table[250]  <= 32'b	00001001100011011101101011101101	;
		random_num_table[251]  <= 32'b	00000011100001011000000010000011	;
		random_num_table[252]  <= 32'b	00001000110011011101100000001110	;
		random_num_table[253]  <= 32'b	00000110100111000101010100110100	;
		random_num_table[254]  <= 32'b	00000111110000110010000110110100	;
		random_num_table[255]  <= 32'b	00011001000010110111100101101111	;
	end
endmodule
