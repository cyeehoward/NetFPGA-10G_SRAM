`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:54:44 01/19/2015 
// Design Name: 
// Module Name:    rand_table_6 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module rand_table_6(axi_aclk , axi_aresetn , index_num , rand_out , en);
	input			axi_aclk , axi_aresetn , en;
	input		[7:0]	index_num;
	output		[31:0]	rand_out;

	reg 		[31:0]	random_num_table  [255:0];

	assign rand_out = en?random_num_table[index_num]:32'd0;
	
	always@(posedge axi_aclk)
	begin
		random_num_table[0]  <= 32'b	00001000101111011100110010010011	;
		random_num_table[1]  <= 32'b	00000101100010100100000000101011	;
		random_num_table[2]  <= 32'b	00010100010001000110101101111101	;
		random_num_table[3]  <= 32'b	00010110110000111000100011101000	;
		random_num_table[4]  <= 32'b	00011111101101100000001001110011	;
		random_num_table[5]  <= 32'b	00000011010101010000001110110000	;
		random_num_table[6]  <= 32'b	00000111011000101100001011010001	;
		random_num_table[7]  <= 32'b	00011000010110001111000100010000	;
		random_num_table[8]  <= 32'b	00011110100101100001011001011001	;
		random_num_table[9]  <= 32'b	00010100110111101100100010110110	;
		random_num_table[10]  <= 32'b	00001010011010110100000010111111	;
		random_num_table[11]  <= 32'b	00000111010000111010111100011101	;
		random_num_table[12]  <= 32'b	00010101101000000111101110111110	;
		random_num_table[13]  <= 32'b	00000111001000011111101010010110	;
		random_num_table[14]  <= 32'b	00000101110100101101000110110100	;
		random_num_table[15]  <= 32'b	00000000110110100101000101000101	;
		random_num_table[16]  <= 32'b	00001111000011010110010110100010	;
		random_num_table[17]  <= 32'b	00010010100011000100100101110111	;
		random_num_table[18]  <= 32'b	00010100100011110011100110100011	;
		random_num_table[19]  <= 32'b	00001110110111001011001010110001	;
		random_num_table[20]  <= 32'b	00001110101111000000100011111110	;
		random_num_table[21]  <= 32'b	00010100010000111000101100111100	;
		random_num_table[22]  <= 32'b	00010100010011111010011111010111	;
		random_num_table[23]  <= 32'b	00001011101010111010110000101110	;
		random_num_table[24]  <= 32'b	00010000100011000000111110001011	;
		random_num_table[25]  <= 32'b	00000111101001011111000011111100	;
		random_num_table[26]  <= 32'b	00010110000001111010000111010001	;
		random_num_table[27]  <= 32'b	00001000001010000110110001100011	;
		random_num_table[28]  <= 32'b	00010010110101100101001111011111	;
		random_num_table[29]  <= 32'b	00000111010100101011110000001111	;
		random_num_table[30]  <= 32'b	00000111110000101111000101101101	;
		random_num_table[31]  <= 32'b	00001100110101100010101100110010	;
		random_num_table[32]  <= 32'b	00000110010001001111010011110010	;
		random_num_table[33]  <= 32'b	00000010100100010100111000110011	;
		random_num_table[34]  <= 32'b	00010111101111011011001101100111	;
		random_num_table[35]  <= 32'b	00001101111001011111011110000110	;
		random_num_table[36]  <= 32'b	00010000010100100101111101000011	;
		random_num_table[37]  <= 32'b	00010000110011101100111010111000	;
		random_num_table[38]  <= 32'b	00010010010101001001011001100001	;
		random_num_table[39]  <= 32'b	00001100101001110100010111101001	;
		random_num_table[40]  <= 32'b	00000101101010111011100100111100	;
		random_num_table[41]  <= 32'b	00001101110101000100011001111010	;
		random_num_table[42]  <= 32'b	00001000110011100100011001011010	;
		random_num_table[43]  <= 32'b	00000110110101110101110001011010	;
		random_num_table[44]  <= 32'b	00010110101101110011110111111100	;
		random_num_table[45]  <= 32'b	00000101100110100000111011001010	;
		random_num_table[46]  <= 32'b	00011111011111010110001010100100	;
		random_num_table[47]  <= 32'b	00011111010110001111100001110100	;
		random_num_table[48]  <= 32'b	00010101110100001101001011010011	;
		random_num_table[49]  <= 32'b	00001100111100001010000110000010	;
		random_num_table[50]  <= 32'b	00001011100101010011100101011111	;
		random_num_table[51]  <= 32'b	00010011010010001001111000011011	;
		random_num_table[52]  <= 32'b	00001011011000010110111011001111	;
		random_num_table[53]  <= 32'b	00001001100001101001101000001111	;
		random_num_table[54]  <= 32'b	00000011110110100100100001001101	;
		random_num_table[55]  <= 32'b	00010001001100100001001011101011	;
		random_num_table[56]  <= 32'b	00000011000000011011011100100011	;
		random_num_table[57]  <= 32'b	00001000100011101100111100111101	;
		random_num_table[58]  <= 32'b	00001010111111100010111101011011	;
		random_num_table[59]  <= 32'b	00010100011110100110001100001010	;
		random_num_table[60]  <= 32'b	00000000100101000011101111110110	;
		random_num_table[61]  <= 32'b	00011010101001011000101000011111	;
		random_num_table[62]  <= 32'b	00001100110100011101100110001101	;
		random_num_table[63]  <= 32'b	00000111011001101010010001010100	;
		random_num_table[64]  <= 32'b	00011001000011011110101001001111	;
		random_num_table[65]  <= 32'b	00011000000011101100110111000001	;
		random_num_table[66]  <= 32'b	00011100110110010110010100101001	;
		random_num_table[67]  <= 32'b	00000111100100100111111011000100	;
		random_num_table[68]  <= 32'b	00001000101101001110011010011101	;
		random_num_table[69]  <= 32'b	00011011111101001101100110101100	;
		random_num_table[70]  <= 32'b	00000110001110100001110111011010	;
		random_num_table[71]  <= 32'b	00010110100111001100010110110110	;
		random_num_table[72]  <= 32'b	00011001011101100101111111110101	;
		random_num_table[73]  <= 32'b	00001111011000010111110000001101	;
		random_num_table[74]  <= 32'b	00000100011001011111100001010011	;
		random_num_table[75]  <= 32'b	00011101111001000101010001000110	;
		random_num_table[76]  <= 32'b	00011111101011001010001101010011	;
		random_num_table[77]  <= 32'b	00001001100001101001111010110110	;
		random_num_table[78]  <= 32'b	00010110111010011011001000000001	;
		random_num_table[79]  <= 32'b	00000110000010010110101100100000	;
		random_num_table[80]  <= 32'b	00001011011001110110100111011101	;
		random_num_table[81]  <= 32'b	00000101110011011011011000111000	;
		random_num_table[82]  <= 32'b	00000101010011000101001011011011	;
		random_num_table[83]  <= 32'b	00010100001111111011000100100111	;
		random_num_table[84]  <= 32'b	00000010101100101011000111101000	;
		random_num_table[85]  <= 32'b	00011100101100010010001011011011	;
		random_num_table[86]  <= 32'b	00010111110110110010000011110011	;
		random_num_table[87]  <= 32'b	00011010110010001111100000101100	;
		random_num_table[88]  <= 32'b	00011001100110010000001010101101	;
		random_num_table[89]  <= 32'b	00011001011110000101101111110111	;
		random_num_table[90]  <= 32'b	00001001001001011111111101110110	;
		random_num_table[91]  <= 32'b	00010000100000010111011100100101	;
		random_num_table[92]  <= 32'b	00000111110111011100100000100100	;
		random_num_table[93]  <= 32'b	00010100000001111011100001101101	;
		random_num_table[94]  <= 32'b	00010111010110110100000010100100	;
		random_num_table[95]  <= 32'b	00000001111101011011101001000010	;
		random_num_table[96]  <= 32'b	00010001010101110110100001000010	;
		random_num_table[97]  <= 32'b	00001100001110000100110011101000	;
		random_num_table[98]  <= 32'b	00010110011001000100000001110000	;
		random_num_table[99]  <= 32'b	00001010011101000000010110101010	;
		random_num_table[100]  <= 32'b	00010111010011000100110110110011	;
		random_num_table[101]  <= 32'b	00010010110100001001101001000011	;
		random_num_table[102]  <= 32'b	00000010111111100000101101011010	;
		random_num_table[103]  <= 32'b	00010110011111100011111001101011	;
		random_num_table[104]  <= 32'b	00000000010001011100100101111000	;
		random_num_table[105]  <= 32'b	00001110110101010010001000101101	;
		random_num_table[106]  <= 32'b	00000111000110110010011100100111	;
		random_num_table[107]  <= 32'b	00000100100011000110101011100010	;
		random_num_table[108]  <= 32'b	00011000000000100110110110001000	;
		random_num_table[109]  <= 32'b	00010111000100100111011111110010	;
		random_num_table[110]  <= 32'b	00001110100111111100100000111011	;
		random_num_table[111]  <= 32'b	00011100001000111101110000101101	;
		random_num_table[112]  <= 32'b	00000110101100110110101010111110	;
		random_num_table[113]  <= 32'b	00000000100101000010100001011100	;
		random_num_table[114]  <= 32'b	00011001101001010100101000001110	;
		random_num_table[115]  <= 32'b	00010101011010010010101110010010	;
		random_num_table[116]  <= 32'b	00000010100101110100011010100100	;
		random_num_table[117]  <= 32'b	00000000100010011011101000100101	;
		random_num_table[118]  <= 32'b	00010101011110111101100000010100	;
		random_num_table[119]  <= 32'b	00010010100100011101110100101001	;
		random_num_table[120]  <= 32'b	00010000001111011101111101011011	;
		random_num_table[121]  <= 32'b	00010010111001001011010010111001	;
		random_num_table[122]  <= 32'b	00001100110000101111000111010100	;
		random_num_table[123]  <= 32'b	00010001000000001111011000100100	;
		random_num_table[124]  <= 32'b	00010101000000011100100110101010	;
		random_num_table[125]  <= 32'b	00000001100110001000101101001100	;
		random_num_table[126]  <= 32'b	00010100000010011011001010010001	;
		random_num_table[127]  <= 32'b	00001100010101011111101010001000	;
		random_num_table[128]  <= 32'b	00000111100011110001010000111010	;
		random_num_table[129]  <= 32'b	00000010110110101110000100100110	;
		random_num_table[130]  <= 32'b	00010111000100111001010100111100	;
		random_num_table[131]  <= 32'b	00001111111011100000011100111011	;
		random_num_table[132]  <= 32'b	00011000100110101000101011000000	;
		random_num_table[133]  <= 32'b	00000110000111000010111011001101	;
		random_num_table[134]  <= 32'b	00010010010000110010111111001001	;
		random_num_table[135]  <= 32'b	00011000101000110001110110000100	;
		random_num_table[136]  <= 32'b	00001100011100000000001111110111	;
		random_num_table[137]  <= 32'b	00011101001110101011100111000101	;
		random_num_table[138]  <= 32'b	00000101110011111111010010000101	;
		random_num_table[139]  <= 32'b	00011101101100001110011111000010	;
		random_num_table[140]  <= 32'b	00001001100110000000010101011100	;
		random_num_table[141]  <= 32'b	00011100011011011101111000011110	;
		random_num_table[142]  <= 32'b	00011011110010100110010100011011	;
		random_num_table[143]  <= 32'b	00001000010100001010000011101010	;
		random_num_table[144]  <= 32'b	00011111100001000101010101000001	;
		random_num_table[145]  <= 32'b	00011010111111000101010101101001	;
		random_num_table[146]  <= 32'b	00011000011011111011100110110101	;
		random_num_table[147]  <= 32'b	00011101000101110010100011010001	;
		random_num_table[148]  <= 32'b	00000110110000001011011111100001	;
		random_num_table[149]  <= 32'b	00000110101011010000100111010110	;
		random_num_table[150]  <= 32'b	00010001110100111111101111101100	;
		random_num_table[151]  <= 32'b	00000101111111010011010001001010	;
		random_num_table[152]  <= 32'b	00010000101100110001010000110111	;
		random_num_table[153]  <= 32'b	00011000001011110100011110010011	;
		random_num_table[154]  <= 32'b	00000111010001110000100011010010	;
		random_num_table[155]  <= 32'b	00001011100110110100111111111101	;
		random_num_table[156]  <= 32'b	00001010001110010101010010001000	;
		random_num_table[157]  <= 32'b	00011010000010011011010001101100	;
		random_num_table[158]  <= 32'b	00001001100101010001101010111100	;
		random_num_table[159]  <= 32'b	00011110011011000111111101001110	;
		random_num_table[160]  <= 32'b	00010001110110101000101111100010	;
		random_num_table[161]  <= 32'b	00001100100100011000010011101001	;
		random_num_table[162]  <= 32'b	00001010111101000011000010011101	;
		random_num_table[163]  <= 32'b	00001111110101111111010110001110	;
		random_num_table[164]  <= 32'b	00011010000000001100000000011010	;
		random_num_table[165]  <= 32'b	00000111011111111010111001010000	;
		random_num_table[166]  <= 32'b	00000110100001000000100100111010	;
		random_num_table[167]  <= 32'b	00000110011100111000000100010001	;
		random_num_table[168]  <= 32'b	00010000111011101111101101000010	;
		random_num_table[169]  <= 32'b	00011111100101000111110101111000	;
		random_num_table[170]  <= 32'b	00000001111011101111001111111111	;
		random_num_table[171]  <= 32'b	00001110100101001111101011111111	;
		random_num_table[172]  <= 32'b	00010001001100110000011010001000	;
		random_num_table[173]  <= 32'b	00000010000010010001100000100111	;
		random_num_table[174]  <= 32'b	00011110001000000000010111011011	;
		random_num_table[175]  <= 32'b	00000010010010110111011110010111	;
		random_num_table[176]  <= 32'b	00000011100011001000101111101011	;
		random_num_table[177]  <= 32'b	00011100010100010111100010000101	;
		random_num_table[178]  <= 32'b	00010001011010000110000110101011	;
		random_num_table[179]  <= 32'b	00011000101001110111011100111011	;
		random_num_table[180]  <= 32'b	00011010111001010011010111000111	;
		random_num_table[181]  <= 32'b	00010010101110100000110011001110	;
		random_num_table[182]  <= 32'b	00001001010100110100101010101011	;
		random_num_table[183]  <= 32'b	00010000111011110111111011100110	;
		random_num_table[184]  <= 32'b	00010001110001010011011110000101	;
		random_num_table[185]  <= 32'b	00000011001110001101000011111011	;
		random_num_table[186]  <= 32'b	00001111101001011001001100100000	;
		random_num_table[187]  <= 32'b	00010011111111111000100001101111	;
		random_num_table[188]  <= 32'b	00000000110001000001010010011001	;
		random_num_table[189]  <= 32'b	00000110001111100010010110001001	;
		random_num_table[190]  <= 32'b	00001101011110100000000110111110	;
		random_num_table[191]  <= 32'b	00010001010101010101100101100111	;
		random_num_table[192]  <= 32'b	00010001101110100000101111100101	;
		random_num_table[193]  <= 32'b	00010000110001110100011110010100	;
		random_num_table[194]  <= 32'b	00001001100011000111000011000010	;
		random_num_table[195]  <= 32'b	00001101010110011111110111011101	;
		random_num_table[196]  <= 32'b	00000111101011010110011010010001	;
		random_num_table[197]  <= 32'b	00000101110010011010101111001001	;
		random_num_table[198]  <= 32'b	00001111000001110111100100000000	;
		random_num_table[199]  <= 32'b	00000001000100100001000000011000	;
		random_num_table[200]  <= 32'b	00010101001110010111010111110110	;
		random_num_table[201]  <= 32'b	00001011101111001001110010100001	;
		random_num_table[202]  <= 32'b	00000010110111101101010000101011	;
		random_num_table[203]  <= 32'b	00000101101010100011101010101000	;
		random_num_table[204]  <= 32'b	00011000001010000010101010010100	;
		random_num_table[205]  <= 32'b	00001001100011010000000101111110	;
		random_num_table[206]  <= 32'b	00001101110001010001001000111010	;
		random_num_table[207]  <= 32'b	00001010111111101011101100111101	;
		random_num_table[208]  <= 32'b	00001100000101011000011110000011	;
		random_num_table[209]  <= 32'b	00000000010101110000010001010100	;
		random_num_table[210]  <= 32'b	00011111000110111110110010001001	;
		random_num_table[211]  <= 32'b	00000110111100101111100000000010	;
		random_num_table[212]  <= 32'b	00000010100101011111010110011001	;
		random_num_table[213]  <= 32'b	00010110000111101110011011110111	;
		random_num_table[214]  <= 32'b	00000101110011111100101100100100	;
		random_num_table[215]  <= 32'b	00001000101111010110000011100000	;
		random_num_table[216]  <= 32'b	00000000101110010000010010000001	;
		random_num_table[217]  <= 32'b	00011111010100011010110010011001	;
		random_num_table[218]  <= 32'b	00011110110010100101001001101110	;
		random_num_table[219]  <= 32'b	00010011001100001000011011110000	;
		random_num_table[220]  <= 32'b	00011001011101110101001100100001	;
		random_num_table[221]  <= 32'b	00001001011010000101110110110001	;
		random_num_table[222]  <= 32'b	00010110011010111111100111011001	;
		random_num_table[223]  <= 32'b	00000011010010000000111001100010	;
		random_num_table[224]  <= 32'b	00000011111010000011101000100110	;
		random_num_table[225]  <= 32'b	00001110111100100110110010010010	;
		random_num_table[226]  <= 32'b	00001101000101101011101011110010	;
		random_num_table[227]  <= 32'b	00000000110000001011101001110101	;
		random_num_table[228]  <= 32'b	00000001101000000011111101000110	;
		random_num_table[229]  <= 32'b	00000110100110000110101011111110	;
		random_num_table[230]  <= 32'b	00000110010001010100111111110001	;
		random_num_table[231]  <= 32'b	00010000001110111110100101110111	;
		random_num_table[232]  <= 32'b	00010010111101100100111001101010	;
		random_num_table[233]  <= 32'b	00000111111101110100101001001111	;
		random_num_table[234]  <= 32'b	00001100110101100001000111000010	;
		random_num_table[235]  <= 32'b	00000110111101011100111110100100	;
		random_num_table[236]  <= 32'b	00000001001011100110010011001110	;
		random_num_table[237]  <= 32'b	00001100010001011100110100010100	;
		random_num_table[238]  <= 32'b	00010010111111000001011111001101	;
		random_num_table[239]  <= 32'b	00000010110000101110101000000010	;
		random_num_table[240]  <= 32'b	00000100011100000000111111010001	;
		random_num_table[241]  <= 32'b	00010011100111111010111010011100	;
		random_num_table[242]  <= 32'b	00001110101011101100001101000001	;
		random_num_table[243]  <= 32'b	00000011000101110010111111000011	;
		random_num_table[244]  <= 32'b	00011010110110000110100001001010	;
		random_num_table[245]  <= 32'b	00011111001010101110111100110100	;
		random_num_table[246]  <= 32'b	00000100001110111111010000000101	;
		random_num_table[247]  <= 32'b	00010010111001100101110110111101	;
		random_num_table[248]  <= 32'b	00000001111011101011001000100100	;
		random_num_table[249]  <= 32'b	00000101100111000000100110101010	;
		random_num_table[250]  <= 32'b	00000101000010111110000101010111	;
		random_num_table[251]  <= 32'b	00001100101001000110010100001111	;
		random_num_table[252]  <= 32'b	00000011101101000000111000011001	;
		random_num_table[253]  <= 32'b	00000101111011000000111011110110	;
		random_num_table[254]  <= 32'b	00000100001010011010010111011010	;
		random_num_table[255]  <= 32'b	00001110110011101111111100101100	;			
	end
endmodule
