`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:54:50 01/19/2015 
// Design Name: 
// Module Name:    rand_table_7 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module rand_table_12(axi_aclk , axi_aresetn , index_num , rand_out , en);
	input			axi_aclk , axi_aresetn , en;
	input		[7:0]	index_num;
	output		[31:0]	rand_out;

	reg 		[31:0]	random_num_table  [255:0];

	assign rand_out = en?random_num_table[index_num]:32'd0;
	
	always@(posedge axi_aclk)
	begin
		random_num_table[0]  <= 32'b	00010111110111111001010001010100	;
		random_num_table[1]  <= 32'b	00000001001000101111011010010110	;
		random_num_table[2]  <= 32'b	00011111000011100100101010100100	;
		random_num_table[3]  <= 32'b	00000101110111100101001110011001	;
		random_num_table[4]  <= 32'b	00011001000110101100011001001100	;
		random_num_table[5]  <= 32'b	00010010010111001011011110001001	;
		random_num_table[6]  <= 32'b	00000100110100001011001100111010	;
		random_num_table[7]  <= 32'b	00001101001010101010011100100001	;
		random_num_table[8]  <= 32'b	00001100001110110100101001111011	;
		random_num_table[9]  <= 32'b	00001100011011010011001100100110	;
		random_num_table[10]  <= 32'b	00010011001110111110110110100011	;
		random_num_table[11]  <= 32'b	00001000001011111000100101000010	;
		random_num_table[12]  <= 32'b	00010001000010110110110110011100	;
		random_num_table[13]  <= 32'b	00001001110011000001110000010101	;
		random_num_table[14]  <= 32'b	00010111010000100110000010011011	;
		random_num_table[15]  <= 32'b	00011111101000111011111011010001	;
		random_num_table[16]  <= 32'b	00001001100011010010110010101110	;
		random_num_table[17]  <= 32'b	00000101000101111111010010011001	;
		random_num_table[18]  <= 32'b	00000101001111010110001111100010	;
		random_num_table[19]  <= 32'b	00011111011110111011110111101011	;
		random_num_table[20]  <= 32'b	00000101000111111001100011111001	;
		random_num_table[21]  <= 32'b	00001001010101110001000111111111	;
		random_num_table[22]  <= 32'b	00001000100010001111010011100100	;
		random_num_table[23]  <= 32'b	00010000000100100100010011001000	;
		random_num_table[24]  <= 32'b	00010000001110010100010000110101	;
		random_num_table[25]  <= 32'b	00000110110001001100111000100010	;
		random_num_table[26]  <= 32'b	00011100110001100010000011100001	;
		random_num_table[27]  <= 32'b	00000001011110000000111111011001	;
		random_num_table[28]  <= 32'b	00001001101010100111100000010010	;
		random_num_table[29]  <= 32'b	00001010111001110111110111000110	;
		random_num_table[30]  <= 32'b	00010111101100100111001010010100	;
		random_num_table[31]  <= 32'b	00010010001000010001000000101101	;
		random_num_table[32]  <= 32'b	00000000111110011100111001101000	;
		random_num_table[33]  <= 32'b	00001011100101001111100110011001	;
		random_num_table[34]  <= 32'b	00010101000111101001000110010011	;
		random_num_table[35]  <= 32'b	00001110001100011000010110110011	;
		random_num_table[36]  <= 32'b	00011101101100110000101100100010	;
		random_num_table[37]  <= 32'b	00000000100100000010110101110011	;
		random_num_table[38]  <= 32'b	00010001101000000010111101010010	;
		random_num_table[39]  <= 32'b	00001001011111101111000100001110	;
		random_num_table[40]  <= 32'b	00010111011111011100110111101001	;
		random_num_table[41]  <= 32'b	00000111111000010110100011010111	;
		random_num_table[42]  <= 32'b	00010001100001111011101100010011	;
		random_num_table[43]  <= 32'b	00000001000000001110001000001111	;
		random_num_table[44]  <= 32'b	00010011011101001011100110111000	;
		random_num_table[45]  <= 32'b	00000110010111000110001110000011	;
		random_num_table[46]  <= 32'b	00000101010110100001010010110101	;
		random_num_table[47]  <= 32'b	00001011010111001001011011000010	;
		random_num_table[48]  <= 32'b	00011010110011110111100111010010	;
		random_num_table[49]  <= 32'b	00010100000110101000110101001001	;
		random_num_table[50]  <= 32'b	00010100001011110011101001010101	;
		random_num_table[51]  <= 32'b	00000000101000110000000011110101	;
		random_num_table[52]  <= 32'b	00011000010100010001011100011010	;
		random_num_table[53]  <= 32'b	00000001010111101110110000001010	;
		random_num_table[54]  <= 32'b	00011101100111000101110110010011	;
		random_num_table[55]  <= 32'b	00001101001100000010000101011100	;
		random_num_table[56]  <= 32'b	00001111000100110000010110111110	;
		random_num_table[57]  <= 32'b	00000100011000010010010001010100	;
		random_num_table[58]  <= 32'b	00001010001011000011111111111001	;
		random_num_table[59]  <= 32'b	00011100010001101001010100100101	;
		random_num_table[60]  <= 32'b	00000100100101001100001101010110	;
		random_num_table[61]  <= 32'b	00011001000100100000110011101110	;
		random_num_table[62]  <= 32'b	00001000000011100111110100011000	;
		random_num_table[63]  <= 32'b	00000010110001010000001000011100	;
		random_num_table[64]  <= 32'b	00001001110010000001110101001001	;
		random_num_table[65]  <= 32'b	00010110011100101110101110010101	;
		random_num_table[66]  <= 32'b	00010100110100101101000011011010	;
		random_num_table[67]  <= 32'b	00011111111101011110010010101000	;
		random_num_table[68]  <= 32'b	00011111011010001100110100100000	;
		random_num_table[69]  <= 32'b	00001010100000011101100101101000	;
		random_num_table[70]  <= 32'b	00001010001101101111001010111000	;
		random_num_table[71]  <= 32'b	00000100011010111101100000010000	;
		random_num_table[72]  <= 32'b	00010110011001101001000000011011	;
		random_num_table[73]  <= 32'b	00010111001011001111111110000111	;
		random_num_table[74]  <= 32'b	00011100100011101011010101010111	;
		random_num_table[75]  <= 32'b	00010110010110000001001001000101	;
		random_num_table[76]  <= 32'b	00000010100110011110101110010111	;
		random_num_table[77]  <= 32'b	00001011011100011001011100000011	;
		random_num_table[78]  <= 32'b	00011100101000111001010111001010	;
		random_num_table[79]  <= 32'b	00011110101111111110101101001010	;
		random_num_table[80]  <= 32'b	00010110001010011011000110101110	;
		random_num_table[81]  <= 32'b	00010111011001010010111000001101	;
		random_num_table[82]  <= 32'b	00001111110110100101100000001001	;
		random_num_table[83]  <= 32'b	00010100001011100001010101111000	;
		random_num_table[84]  <= 32'b	00001100011010011000011011010111	;
		random_num_table[85]  <= 32'b	00010001001110011110001111110011	;
		random_num_table[86]  <= 32'b	00000101111110001100010011100011	;
		random_num_table[87]  <= 32'b	00010000101101111000000100111111	;
		random_num_table[88]  <= 32'b	00001101111010110111101100000000	;
		random_num_table[89]  <= 32'b	00000110011000011101110001001000	;
		random_num_table[90]  <= 32'b	00000110111011000001100110110110	;
		random_num_table[91]  <= 32'b	00001011000010100111000101111100	;
		random_num_table[92]  <= 32'b	00000011100011101000000101011110	;
		random_num_table[93]  <= 32'b	00010111110000111101111110111011	;
		random_num_table[94]  <= 32'b	00001000101101111101111011110001	;
		random_num_table[95]  <= 32'b	00000111000111110111001001000001	;
		random_num_table[96]  <= 32'b	00001101101000010110101111011001	;
		random_num_table[97]  <= 32'b	00010101100110111000110111101100	;
		random_num_table[98]  <= 32'b	00010010011100000110111011101100	;
		random_num_table[99]  <= 32'b	00000111011110101010100010011101	;
		random_num_table[100]  <= 32'b	00011001000100101011111000001101	;
		random_num_table[101]  <= 32'b	00000111011011111101101111100010	;
		random_num_table[102]  <= 32'b	00011010111101010101010100101110	;
		random_num_table[103]  <= 32'b	00001111100001001011011110001110	;
		random_num_table[104]  <= 32'b	00000000001011100110001000000000	;
		random_num_table[105]  <= 32'b	00000001010111000111111001001010	;
		random_num_table[106]  <= 32'b	00011011100101011100000100111011	;
		random_num_table[107]  <= 32'b	00001111001001001010101011100001	;
		random_num_table[108]  <= 32'b	00011000001011111111100100011101	;
		random_num_table[109]  <= 32'b	00010110101011001101110111011100	;
		random_num_table[110]  <= 32'b	00001000011101000100111100010111	;
		random_num_table[111]  <= 32'b	00000101110000001110000111001101	;
		random_num_table[112]  <= 32'b	00010000000111001101101010111000	;
		random_num_table[113]  <= 32'b	00000101001011101101011000001100	;
		random_num_table[114]  <= 32'b	00011000000000101101101010111101	;
		random_num_table[115]  <= 32'b	00011101011100101101100100000100	;
		random_num_table[116]  <= 32'b	00001010011000110101101001000000	;
		random_num_table[117]  <= 32'b	00010010101011111001110001111100	;
		random_num_table[118]  <= 32'b	00010110111001010010111110111010	;
		random_num_table[119]  <= 32'b	00010011000001000000110110110010	;
		random_num_table[120]  <= 32'b	00010110011101101011111010011011	;
		random_num_table[121]  <= 32'b	00010110010101001110001101100010	;
		random_num_table[122]  <= 32'b	00011111100001000101001110100001	;
		random_num_table[123]  <= 32'b	00001001101111111011111001011110	;
		random_num_table[124]  <= 32'b	00011010000110011011010010100010	;
		random_num_table[125]  <= 32'b	00010101001101100111010111101100	;
		random_num_table[126]  <= 32'b	00011011010100110000100101110110	;
		random_num_table[127]  <= 32'b	00011110011011110110011101011111	;
		random_num_table[128]  <= 32'b	00011010010100001111001101001110	;
		random_num_table[129]  <= 32'b	00011100111001101110001010100111	;
		random_num_table[130]  <= 32'b	00010000110001001101000011000001	;
		random_num_table[131]  <= 32'b	00001010000101110011111001001111	;
		random_num_table[132]  <= 32'b	00000111110001000111101001100000	;
		random_num_table[133]  <= 32'b	00010100100000010101011011001000	;
		random_num_table[134]  <= 32'b	00000001011111011001011000010010	;
		random_num_table[135]  <= 32'b	00011011011000111110111010011011	;
		random_num_table[136]  <= 32'b	00011010111011101001100010000100	;
		random_num_table[137]  <= 32'b	00010100011111010110010011111001	;
		random_num_table[138]  <= 32'b	00011110101111110000000001010000	;
		random_num_table[139]  <= 32'b	00011111100101101000101000010010	;
		random_num_table[140]  <= 32'b	00001010111110010011000100110100	;
		random_num_table[141]  <= 32'b	00000000000110010110111011000010	;
		random_num_table[142]  <= 32'b	00001000000110100111101110010110	;
		random_num_table[143]  <= 32'b	00011000011011101000101011101101	;
		random_num_table[144]  <= 32'b	00000011000100110001011010000110	;
		random_num_table[145]  <= 32'b	00011000001110111010001010010100	;
		random_num_table[146]  <= 32'b	00010011001101101001111100111010	;
		random_num_table[147]  <= 32'b	00001100100101110011101000011001	;
		random_num_table[148]  <= 32'b	00011011011100100100110011011001	;
		random_num_table[149]  <= 32'b	00010101101000010111101101010000	;
		random_num_table[150]  <= 32'b	00000101000101101101000011000100	;
		random_num_table[151]  <= 32'b	00000100101000000101101110100011	;
		random_num_table[152]  <= 32'b	00011000101110100111001101101111	;
		random_num_table[153]  <= 32'b	00010000010111101110010001111011	;
		random_num_table[154]  <= 32'b	00011100001000001100111001111001	;
		random_num_table[155]  <= 32'b	00010101111111101000111111101011	;
		random_num_table[156]  <= 32'b	00011001000100001000010000101110	;
		random_num_table[157]  <= 32'b	00011110111000111010100000101101	;
		random_num_table[158]  <= 32'b	00010011011111100010001001001001	;
		random_num_table[159]  <= 32'b	00001100011111000101101111011010	;
		random_num_table[160]  <= 32'b	00010110000011101011110011100100	;
		random_num_table[161]  <= 32'b	00011010101010010000011111111001	;
		random_num_table[162]  <= 32'b	00010001110111111101100101011110	;
		random_num_table[163]  <= 32'b	00001101111110111011100010010110	;
		random_num_table[164]  <= 32'b	00000001010010100110011001010001	;
		random_num_table[165]  <= 32'b	00011110011110111110100100001111	;
		random_num_table[166]  <= 32'b	00000101000100110011100001101011	;
		random_num_table[167]  <= 32'b	00011111010110101010111101011011	;
		random_num_table[168]  <= 32'b	00001011101011011110111100010001	;
		random_num_table[169]  <= 32'b	00001001110001010110101100111000	;
		random_num_table[170]  <= 32'b	00011111101010100000011101111011	;
		random_num_table[171]  <= 32'b	00010010001100100100111011110011	;
		random_num_table[172]  <= 32'b	00010101000110101001011110110010	;
		random_num_table[173]  <= 32'b	00000011011000000111010110010000	;
		random_num_table[174]  <= 32'b	00000110000111000111000010011001	;
		random_num_table[175]  <= 32'b	00000110100011010011111111000110	;
		random_num_table[176]  <= 32'b	00010010101010110101001110011100	;
		random_num_table[177]  <= 32'b	00000101010110010110100000001010	;
		random_num_table[178]  <= 32'b	00010011010101011101100111111101	;
		random_num_table[179]  <= 32'b	00001000010011111001110011100111	;
		random_num_table[180]  <= 32'b	00000001010010111110101001111010	;
		random_num_table[181]  <= 32'b	00001100101001000000011100001010	;
		random_num_table[182]  <= 32'b	00010001111011001111010000010110	;
		random_num_table[183]  <= 32'b	00001000011000101011001011011001	;
		random_num_table[184]  <= 32'b	00001100011111010101111001101101	;
		random_num_table[185]  <= 32'b	00011101011101011001010101011111	;
		random_num_table[186]  <= 32'b	00011110100111010111011110001000	;
		random_num_table[187]  <= 32'b	00001101010011101010001110001111	;
		random_num_table[188]  <= 32'b	00000111000010100011001010111011	;
		random_num_table[189]  <= 32'b	00001100000000110010100101000010	;
		random_num_table[190]  <= 32'b	00001101110101011000001111011100	;
		random_num_table[191]  <= 32'b	00010000001001001010110010100000	;
		random_num_table[192]  <= 32'b	00010010001111011101001101111010	;
		random_num_table[193]  <= 32'b	00000000101011100100110111110001	;
		random_num_table[194]  <= 32'b	00001110001011000000011100010111	;
		random_num_table[195]  <= 32'b	00011101000000110111101100101001	;
		random_num_table[196]  <= 32'b	00010010011100010100000101100100	;
		random_num_table[197]  <= 32'b	00011111111110110010011101111110	;
		random_num_table[198]  <= 32'b	00001100011101111110010010111101	;
		random_num_table[199]  <= 32'b	00001001110101000101011001001101	;
		random_num_table[200]  <= 32'b	00001000111011000101000101110010	;
		random_num_table[201]  <= 32'b	00011101010011011011101001001000	;
		random_num_table[202]  <= 32'b	00010001001010100011101000011100	;
		random_num_table[203]  <= 32'b	00001010101111111111011001110101	;
		random_num_table[204]  <= 32'b	00010001100010111010011011000001	;
		random_num_table[205]  <= 32'b	00010101100000001101010100110101	;
		random_num_table[206]  <= 32'b	00010000011101110111000011011011	;
		random_num_table[207]  <= 32'b	00000101110100000010101101000101	;
		random_num_table[208]  <= 32'b	00011110110101101011000110010011	;
		random_num_table[209]  <= 32'b	00011111001100111111111010001000	;
		random_num_table[210]  <= 32'b	00010100001101110111101100101011	;
		random_num_table[211]  <= 32'b	00011001000001001011000010110001	;
		random_num_table[212]  <= 32'b	00000001001000110110100000110000	;
		random_num_table[213]  <= 32'b	00010110101000101000110010101000	;
		random_num_table[214]  <= 32'b	00000110000110101011001101000101	;
		random_num_table[215]  <= 32'b	00010001100011101001111010011100	;
		random_num_table[216]  <= 32'b	00001001011110011101010001001010	;
		random_num_table[217]  <= 32'b	00001010011111010010001011101111	;
		random_num_table[218]  <= 32'b	00011111110011001101010101010000	;
		random_num_table[219]  <= 32'b	00011000001000111000010001110111	;
		random_num_table[220]  <= 32'b	00001000101001110001011001010110	;
		random_num_table[221]  <= 32'b	00001111101101100001001100001011	;
		random_num_table[222]  <= 32'b	00001110100000000011010111111101	;
		random_num_table[223]  <= 32'b	00010110101111110101100110101010	;
		random_num_table[224]  <= 32'b	00011011110011011001100010000110	;
		random_num_table[225]  <= 32'b	00010011000101001100101100010011	;
		random_num_table[226]  <= 32'b	00001110100110100010100001100111	;
		random_num_table[227]  <= 32'b	00000000110000111110000100101010	;
		random_num_table[228]  <= 32'b	00010100101101111010110011110100	;
		random_num_table[229]  <= 32'b	00001010000011010101101011011010	;
		random_num_table[230]  <= 32'b	00001001101010010010011000110110	;
		random_num_table[231]  <= 32'b	00010111101100011011001011000100	;
		random_num_table[232]  <= 32'b	00001010100011111001110101010001	;
		random_num_table[233]  <= 32'b	00000100010110010111011100010011	;
		random_num_table[234]  <= 32'b	00011100001100010010100011011011	;
		random_num_table[235]  <= 32'b	00010110011111010101111011011011	;
		random_num_table[236]  <= 32'b	00001111000110010111111011010100	;
		random_num_table[237]  <= 32'b	00011010101001011101001111100010	;
		random_num_table[238]  <= 32'b	00000110001010011011101101100111	;
		random_num_table[239]  <= 32'b	00001101010001110100000100011100	;
		random_num_table[240]  <= 32'b	00011011011100011111001011110010	;
		random_num_table[241]  <= 32'b	00011001000110110001000000010010	;
		random_num_table[242]  <= 32'b	00010111100111111110011011010101	;
		random_num_table[243]  <= 32'b	00011110100011110110010101000000	;
		random_num_table[244]  <= 32'b	00000010011000110100110011111101	;
		random_num_table[245]  <= 32'b	00001101001101000100010000110010	;
		random_num_table[246]  <= 32'b	00010000101000001111101110011010	;
		random_num_table[247]  <= 32'b	00001110101000100110000100100111	;
		random_num_table[248]  <= 32'b	00001010001010001101010010001111	;
		random_num_table[249]  <= 32'b	00001000001011011100110110100010	;
		random_num_table[250]  <= 32'b	00011100111110110010100001111011	;
		random_num_table[251]  <= 32'b	00000011100101010111101010000000	;
		random_num_table[252]  <= 32'b	00001011100111011001110100111100	;
		random_num_table[253]  <= 32'b	00010101111110001011001100011001	;
		random_num_table[254]  <= 32'b	00010101000001010111111000011011	;
		random_num_table[255]  <= 32'b	00001101000110101101001110111110	;			
	end
endmodule
