`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:54:50 01/19/2015 
// Design Name: 
// Module Name:    rand_table_7 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module rand_table_10(axi_aclk , axi_aresetn , index_num , rand_out , en);
	input			axi_aclk , axi_aresetn , en;
	input		[7:0]	index_num;
	output		[31:0]	rand_out;

	reg 		[31:0]	random_num_table  [255:0];

	assign rand_out = en?random_num_table[index_num]:32'd0;
	
	always@(posedge axi_aclk)
	begin
		random_num_table[0]  <= 32'b	00011011011011101101111101101010	;
		random_num_table[1]  <= 32'b	00010010100001000100001100111111	;
		random_num_table[2]  <= 32'b	00010011010000111001100111110110	;
		random_num_table[3]  <= 32'b	00001011110101010111100100111010	;
		random_num_table[4]  <= 32'b	00011111110000001001001100111010	;
		random_num_table[5]  <= 32'b	00000101010011101111011101101011	;
		random_num_table[6]  <= 32'b	00000100100101000100100101001101	;
		random_num_table[7]  <= 32'b	00001101010011010011110110010010	;
		random_num_table[8]  <= 32'b	00010111000000100000101010000000	;
		random_num_table[9]  <= 32'b	00001100010011101101000100001100	;
		random_num_table[10]  <= 32'b	00011110100111100011110001010110	;
		random_num_table[11]  <= 32'b	00001111000000001101001010000011	;
		random_num_table[12]  <= 32'b	00010001100000010001001011101101	;
		random_num_table[13]  <= 32'b	00000001001111110011010111100011	;
		random_num_table[14]  <= 32'b	00011101110111100100000100100011	;
		random_num_table[15]  <= 32'b	00010100010011110101100111001101	;
		random_num_table[16]  <= 32'b	00011010110010101001110111101010	;
		random_num_table[17]  <= 32'b	00011111000110110100100101110101	;
		random_num_table[18]  <= 32'b	00010101110001010100100000010011	;
		random_num_table[19]  <= 32'b	00000001110100001111111010000110	;
		random_num_table[20]  <= 32'b	00010010111000010000000000101000	;
		random_num_table[21]  <= 32'b	00000010010111101000110001001111	;
		random_num_table[22]  <= 32'b	00000100101010000110011100011010	;
		random_num_table[23]  <= 32'b	00010011000001110000111001001100	;
		random_num_table[24]  <= 32'b	00010011000110110110001000100111	;
		random_num_table[25]  <= 32'b	00001100100010111110011011010010	;
		random_num_table[26]  <= 32'b	00011001000110100010101110010101	;
		random_num_table[27]  <= 32'b	00010000110010100011011111111000	;
		random_num_table[28]  <= 32'b	00011111111001001101100100111010	;
		random_num_table[29]  <= 32'b	00011111101100011011010000111010	;
		random_num_table[30]  <= 32'b	00000001001001101011111101110101	;
		random_num_table[31]  <= 32'b	00000101101000110000110101000111	;
		random_num_table[32]  <= 32'b	00011000101000001011001001110111	;
		random_num_table[33]  <= 32'b	00000011110110110010111111111000	;
		random_num_table[34]  <= 32'b	00010001101101100101100000011101	;
		random_num_table[35]  <= 32'b	00000000101000110100000000011001	;
		random_num_table[36]  <= 32'b	00001011111100101011100101111010	;
		random_num_table[37]  <= 32'b	00011110111000100100100011000111	;
		random_num_table[38]  <= 32'b	00011101100010100101011010010111	;
		random_num_table[39]  <= 32'b	00001100100011100110111000111011	;
		random_num_table[40]  <= 32'b	00000001101001010011010011111110	;
		random_num_table[41]  <= 32'b	00000001101100000011010010100100	;
		random_num_table[42]  <= 32'b	00010000011100010110111000010100	;
		random_num_table[43]  <= 32'b	00001011101111011001001010110001	;
		random_num_table[44]  <= 32'b	00000001010000001000101011010100	;
		random_num_table[45]  <= 32'b	00011000011101001111111010111010	;
		random_num_table[46]  <= 32'b	00010001010001110001011001101000	;
		random_num_table[47]  <= 32'b	00001100111111101000010011000111	;
		random_num_table[48]  <= 32'b	00000100001001010100001001111110	;
		random_num_table[49]  <= 32'b	00001110110010001110111100100110	;
		random_num_table[50]  <= 32'b	00010101101011001110100011111001	;
		random_num_table[51]  <= 32'b	00000100110011011110000100100000	;
		random_num_table[52]  <= 32'b	00011000101010000100001111111110	;
		random_num_table[53]  <= 32'b	00000010011010101101000110001000	;
		random_num_table[54]  <= 32'b	00000011111001011011000001011000	;
		random_num_table[55]  <= 32'b	00000010010100111101100011101010	;
		random_num_table[56]  <= 32'b	00001101100100100001100001000000	;
		random_num_table[57]  <= 32'b	00001100001000011100111001111111	;
		random_num_table[58]  <= 32'b	00001111101000010010000100100011	;
		random_num_table[59]  <= 32'b	00000101000010010110111101001100	;
		random_num_table[60]  <= 32'b	00010100000010000010010100110111	;
		random_num_table[61]  <= 32'b	00011011110100011110000011000010	;
		random_num_table[62]  <= 32'b	00011111011011011111111001110011	;
		random_num_table[63]  <= 32'b	00011000001000000111110001010011	;
		random_num_table[64]  <= 32'b	00001101100010011010011011101100	;
		random_num_table[65]  <= 32'b	00001101001001100110100101110100	;
		random_num_table[66]  <= 32'b	00010100011111000111100100011101	;
		random_num_table[67]  <= 32'b	00010001110001101010101100110100	;
		random_num_table[68]  <= 32'b	00001011001000101100000100101111	;
		random_num_table[69]  <= 32'b	00011111111110111110010100001010	;
		random_num_table[70]  <= 32'b	00011011011011001110110111001111	;
		random_num_table[71]  <= 32'b	00000101011011100001111001001101	;
		random_num_table[72]  <= 32'b	00010000101001001010111001000100	;
		random_num_table[73]  <= 32'b	00011110100000001001101011110001	;
		random_num_table[74]  <= 32'b	00000010101110110101000001111100	;
		random_num_table[75]  <= 32'b	00001011101010000101010010001100	;
		random_num_table[76]  <= 32'b	00010011111001100110110000110101	;
		random_num_table[77]  <= 32'b	00010101111011100001011101011000	;
		random_num_table[78]  <= 32'b	00011011011011100101011111000011	;
		random_num_table[79]  <= 32'b	00000001111001101011000010001100	;
		random_num_table[80]  <= 32'b	00011000110110011100010010000100	;
		random_num_table[81]  <= 32'b	00000001001010000101010111111000	;
		random_num_table[82]  <= 32'b	00000101000000000000101010110100	;
		random_num_table[83]  <= 32'b	00010001110100111110010100100100	;
		random_num_table[84]  <= 32'b	00000100010010000100010100101010	;
		random_num_table[85]  <= 32'b	00001110000110011011111110000111	;
		random_num_table[86]  <= 32'b	00010000110100110011110000100010	;
		random_num_table[87]  <= 32'b	00001111011001010111110111101001	;
		random_num_table[88]  <= 32'b	00000011000111110011101111001110	;
		random_num_table[89]  <= 32'b	00011100011110010111110110110010	;
		random_num_table[90]  <= 32'b	00011000100110111111111011100000	;
		random_num_table[91]  <= 32'b	00010101110100100001001101000101	;
		random_num_table[92]  <= 32'b	00000101101111011011110100000101	;
		random_num_table[93]  <= 32'b	00011100001000100010101011111000	;
		random_num_table[94]  <= 32'b	00010101011100110100010101010101	;
		random_num_table[95]  <= 32'b	00011000101011011110111101100111	;
		random_num_table[96]  <= 32'b	00001111010010000010100011100010	;
		random_num_table[97]  <= 32'b	00001010000011101111110101101001	;
		random_num_table[98]  <= 32'b	00000101111000000010000111001000	;
		random_num_table[99]  <= 32'b	00011011001011011101101110110011	;
		random_num_table[100]  <= 32'b	00001101000001000110110011110011	;
		random_num_table[101]  <= 32'b	00010011110101111001001010010000	;
		random_num_table[102]  <= 32'b	00010011100000011110010110111001	;
		random_num_table[103]  <= 32'b	00000011010111010010100011100110	;
		random_num_table[104]  <= 32'b	00001011101101010110000101000000	;
		random_num_table[105]  <= 32'b	00010101101110011000000000000011	;
		random_num_table[106]  <= 32'b	00001100101111001111000111110100	;
		random_num_table[107]  <= 32'b	00000010100010101100100011011011	;
		random_num_table[108]  <= 32'b	00001110110011100011000001101000	;
		random_num_table[109]  <= 32'b	00010010100111000011100101101011	;
		random_num_table[110]  <= 32'b	00010000110011000010000010110001	;
		random_num_table[111]  <= 32'b	00001101100001110100111100100010	;
		random_num_table[112]  <= 32'b	00010011000110000101101010010100	;
		random_num_table[113]  <= 32'b	00000110001101011011110111000000	;
		random_num_table[114]  <= 32'b	00000000001001100101001010110001	;
		random_num_table[115]  <= 32'b	00000110111101010100001011001001	;
		random_num_table[116]  <= 32'b	00010001100100100110010101010111	;
		random_num_table[117]  <= 32'b	00011111100100111111101000011000	;
		random_num_table[118]  <= 32'b	00000011110101100011110011100010	;
		random_num_table[119]  <= 32'b	00001001100010110001110110100100	;
		random_num_table[120]  <= 32'b	00010001011110000110100111100000	;
		random_num_table[121]  <= 32'b	00000011000111011110101110011011	;
		random_num_table[122]  <= 32'b	00010100110111011001101110010100	;
		random_num_table[123]  <= 32'b	00010100010001100010001111010000	;
		random_num_table[124]  <= 32'b	00010101001111100110111101011111	;
		random_num_table[125]  <= 32'b	00010011011101010111011001000110	;
		random_num_table[126]  <= 32'b	00001111001000111100001100111101	;
		random_num_table[127]  <= 32'b	00001001111111001101010011010101	;
		random_num_table[128]  <= 32'b	00001001011101001010111010100110	;
		random_num_table[129]  <= 32'b	00011110100101101100111011101111	;
		random_num_table[130]  <= 32'b	00010100000011000101011011100110	;
		random_num_table[131]  <= 32'b	00000011000101110001010100011011	;
		random_num_table[132]  <= 32'b	00010111010010101101011011001001	;
		random_num_table[133]  <= 32'b	00010000010001111010010100010101	;
		random_num_table[134]  <= 32'b	00000101011001100011110101100001	;
		random_num_table[135]  <= 32'b	00011101111000001111110101100010	;
		random_num_table[136]  <= 32'b	00011011010010011010011101010111	;
		random_num_table[137]  <= 32'b	00001010000001011101000101001100	;
		random_num_table[138]  <= 32'b	00000100101010111110100000110100	;
		random_num_table[139]  <= 32'b	00001111111011100010010110110011	;
		random_num_table[140]  <= 32'b	00001011101011101001101000101011	;
		random_num_table[141]  <= 32'b	00011000011101101111000010100110	;
		random_num_table[142]  <= 32'b	00010100100011110111001010110100	;
		random_num_table[143]  <= 32'b	00001001100011100001101011010110	;
		random_num_table[144]  <= 32'b	00001110100110101111101100011010	;
		random_num_table[145]  <= 32'b	00010110010111110101100011000011	;
		random_num_table[146]  <= 32'b	00011010110110111011101010100010	;
		random_num_table[147]  <= 32'b	00000110011101011000111101100001	;
		random_num_table[148]  <= 32'b	00000111101011011101001101111000	;
		random_num_table[149]  <= 32'b	00011101011110011110000100011101	;
		random_num_table[150]  <= 32'b	00010011101010101010001111111100	;
		random_num_table[151]  <= 32'b	00010001101001001000111011101110	;
		random_num_table[152]  <= 32'b	00000010111011100110011101111110	;
		random_num_table[153]  <= 32'b	00011000010001111001001101000010	;
		random_num_table[154]  <= 32'b	00010100111011001111110110111110	;
		random_num_table[155]  <= 32'b	00001000101010001101111100010010	;
		random_num_table[156]  <= 32'b	00001011110110010100001101110110	;
		random_num_table[157]  <= 32'b	00011110001001011100010100110011	;
		random_num_table[158]  <= 32'b	00011101010100101001100010010000	;
		random_num_table[159]  <= 32'b	00011100010000010001110010100000	;
		random_num_table[160]  <= 32'b	00011000010110111110011011001010	;
		random_num_table[161]  <= 32'b	00011001011111100110110010101100	;
		random_num_table[162]  <= 32'b	00000111110010000101011011001101	;
		random_num_table[163]  <= 32'b	00011111000111001010000110001101	;
		random_num_table[164]  <= 32'b	00001110001110010111001111100011	;
		random_num_table[165]  <= 32'b	00001101110011101010010011110000	;
		random_num_table[166]  <= 32'b	00010001001110110111011111011100	;
		random_num_table[167]  <= 32'b	00000001100100001111001100111000	;
		random_num_table[168]  <= 32'b	00011011100111011111111110000111	;
		random_num_table[169]  <= 32'b	00001111110111001011101111111101	;
		random_num_table[170]  <= 32'b	00011111101000001000011000100001	;
		random_num_table[171]  <= 32'b	00001101110101001001010000100111	;
		random_num_table[172]  <= 32'b	00010101001111101010000011110011	;
		random_num_table[173]  <= 32'b	00010011010111011010110010100010	;
		random_num_table[174]  <= 32'b	00000000000111110011101101111001	;
		random_num_table[175]  <= 32'b	00011000110100110101000010101010	;
		random_num_table[176]  <= 32'b	00011000100000111000011011110011	;
		random_num_table[177]  <= 32'b	00000011111001000010111111111110	;
		random_num_table[178]  <= 32'b	00011011100111100000001010111010	;
		random_num_table[179]  <= 32'b	00011001010000111010100110010101	;
		random_num_table[180]  <= 32'b	00010011110110100001111111110111	;
		random_num_table[181]  <= 32'b	00011000010001000111001110110100	;
		random_num_table[182]  <= 32'b	00001110100100110010110001101111	;
		random_num_table[183]  <= 32'b	00001011110100001110110111000110	;
		random_num_table[184]  <= 32'b	00000000001111110100010001111111	;
		random_num_table[185]  <= 32'b	00000110101101011001000101010001	;
		random_num_table[186]  <= 32'b	00010110001010100101111100111010	;
		random_num_table[187]  <= 32'b	00011000011000011111000001011001	;
		random_num_table[188]  <= 32'b	00011010001101110101010101111111	;
		random_num_table[189]  <= 32'b	00010000000100101001011000111101	;
		random_num_table[190]  <= 32'b	00001010010001101101010011111101	;
		random_num_table[191]  <= 32'b	00001000010101111001111001000011	;
		random_num_table[192]  <= 32'b	00001011011111111101000110010011	;
		random_num_table[193]  <= 32'b	00001000010111110111111111001000	;
		random_num_table[194]  <= 32'b	00001111001100100101110000111000	;
		random_num_table[195]  <= 32'b	00000111100101111101101000010110	;
		random_num_table[196]  <= 32'b	00000111101000100101110100110000	;
		random_num_table[197]  <= 32'b	00011001100101101100101000110111	;
		random_num_table[198]  <= 32'b	00010111100001111010010111101010	;
		random_num_table[199]  <= 32'b	00011001001100101011100001110010	;
		random_num_table[200]  <= 32'b	00010101111111110010001011100011	;
		random_num_table[201]  <= 32'b	00011111110000001100110110010101	;
		random_num_table[202]  <= 32'b	00000011011001000000000101000100	;
		random_num_table[203]  <= 32'b	00000111110001010110111110111001	;
		random_num_table[204]  <= 32'b	00001011100111101001100010110011	;
		random_num_table[205]  <= 32'b	00010100010101001011110001001110	;
		random_num_table[206]  <= 32'b	00000110010110001000000110011110	;
		random_num_table[207]  <= 32'b	00010110000001110000010100111000	;
		random_num_table[208]  <= 32'b	00010000110101011101001001110100	;
		random_num_table[209]  <= 32'b	00001011011010100010011000101010	;
		random_num_table[210]  <= 32'b	00010000000011000011100001111000	;
		random_num_table[211]  <= 32'b	00000001111100000110100110111000	;
		random_num_table[212]  <= 32'b	00011010100010110010100001110111	;
		random_num_table[213]  <= 32'b	00011110100011110011110001101011	;
		random_num_table[214]  <= 32'b	00000101001100010011101100011101	;
		random_num_table[215]  <= 32'b	00001010110001001011000011110001	;
		random_num_table[216]  <= 32'b	00001011001101000011110100101100	;
		random_num_table[217]  <= 32'b	00011101111100100101010001111100	;
		random_num_table[218]  <= 32'b	00010100111010100110101100100100	;
		random_num_table[219]  <= 32'b	00010001000111101001100011001000	;
		random_num_table[220]  <= 32'b	00010011100000111011000110110011	;
		random_num_table[221]  <= 32'b	00001110010010110101100001000011	;
		random_num_table[222]  <= 32'b	00001011001011110110100110000110	;
		random_num_table[223]  <= 32'b	00001110110111011111010010000110	;
		random_num_table[224]  <= 32'b	00011000000010110101001100111010	;
		random_num_table[225]  <= 32'b	00010011100000100010011100101101	;
		random_num_table[226]  <= 32'b	00001101000100101101001101010101	;
		random_num_table[227]  <= 32'b	00010011001011100101111011100100	;
		random_num_table[228]  <= 32'b	00011111110111111000001000110110	;
		random_num_table[229]  <= 32'b	00011101011010110010010011010100	;
		random_num_table[230]  <= 32'b	00011101100110111010000100101000	;
		random_num_table[231]  <= 32'b	00010001101101010011010101000001	;
		random_num_table[232]  <= 32'b	00000001000110011111101010110010	;
		random_num_table[233]  <= 32'b	00000011101100101111000010111011	;
		random_num_table[234]  <= 32'b	00011101010111110001010101011110	;
		random_num_table[235]  <= 32'b	00011110000000110001110110001110	;
		random_num_table[236]  <= 32'b	00011101111000101110011001000111	;
		random_num_table[237]  <= 32'b	00000100010011010000111011111011	;
		random_num_table[238]  <= 32'b	00011101000000001001001001001011	;
		random_num_table[239]  <= 32'b	00011101001001110100111101011111	;
		random_num_table[240]  <= 32'b	00001011001010100110010100110011	;
		random_num_table[241]  <= 32'b	00010010001011001101001001101001	;
		random_num_table[242]  <= 32'b	00001010010011000110101101100100	;
		random_num_table[243]  <= 32'b	00001101010111001110001100101010	;
		random_num_table[244]  <= 32'b	00001100001001011011110000010000	;
		random_num_table[245]  <= 32'b	00011110101100101011001100011010	;
		random_num_table[246]  <= 32'b	00010111001101000010000000001000	;
		random_num_table[247]  <= 32'b	00000111010001000110000001010100	;
		random_num_table[248]  <= 32'b	00001010001001000011110101101101	;
		random_num_table[249]  <= 32'b	00000101010000011001001110101110	;
		random_num_table[250]  <= 32'b	00001010011110110000111001101010	;
		random_num_table[251]  <= 32'b	00000111010101110101110010111000	;
		random_num_table[252]  <= 32'b	00001100100011100001111011010011	;
		random_num_table[253]  <= 32'b	00010100001010110000101111000110	;
		random_num_table[254]  <= 32'b	00001011010110011110110100010110	;
		random_num_table[255]  <= 32'b	00011001001110110000000100000100	;			
	end
endmodule
