`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:54:50 01/19/2015 
// Design Name: 
// Module Name:    rand_table_7 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module rand_table_8(axi_aclk , axi_aresetn , index_num , rand_out , en);
	input			axi_aclk , axi_aresetn , en;
	input		[7:0]	index_num;
	output		[31:0]	rand_out;

	reg 		[31:0]	random_num_table  [255:0];

	assign rand_out = en?random_num_table[index_num]:32'd0;
	
	always@(posedge axi_aclk)
	begin
		random_num_table[0]  <= 32'b	00001101101110101100010101110010	;
		random_num_table[1]  <= 32'b	00010101001011110110001000110011	;
		random_num_table[2]  <= 32'b	00010011111011001101110100011111	;
		random_num_table[3]  <= 32'b	00011100100011111111100110111001	;
		random_num_table[4]  <= 32'b	00001000110010000001110111001010	;
		random_num_table[5]  <= 32'b	00010101100010100011001000110001	;
		random_num_table[6]  <= 32'b	00000001000101110100001010010001	;
		random_num_table[7]  <= 32'b	00010010011010010100011010000001	;
		random_num_table[8]  <= 32'b	00000001101010100111110110011000	;
		random_num_table[9]  <= 32'b	00001111100011010011101011101100	;
		random_num_table[10]  <= 32'b	00000000100011001010000001011110	;
		random_num_table[11]  <= 32'b	00000100111011100101000101111111	;
		random_num_table[12]  <= 32'b	00001111010000000010001001100000	;
		random_num_table[13]  <= 32'b	00010010001111110110001000101100	;
		random_num_table[14]  <= 32'b	00011010100101110101111110010101	;
		random_num_table[15]  <= 32'b	00011101011000011110010110111100	;
		random_num_table[16]  <= 32'b	00010010100010111100001001111111	;
		random_num_table[17]  <= 32'b	00010000010100010110000010101111	;
		random_num_table[18]  <= 32'b	00001101010000000100000001110111	;
		random_num_table[19]  <= 32'b	00010011111111100011011000010011	;
		random_num_table[20]  <= 32'b	00010101011011010111001111110101	;
		random_num_table[21]  <= 32'b	00001101001000011010111000010010	;
		random_num_table[22]  <= 32'b	00001110101011100111101100001110	;
		random_num_table[23]  <= 32'b	00000010101100111001110100011011	;
		random_num_table[24]  <= 32'b	00010001010110101010000110100010	;
		random_num_table[25]  <= 32'b	00010000000010110001000111000001	;
		random_num_table[26]  <= 32'b	00000100001110010000010000101110	;
		random_num_table[27]  <= 32'b	00001000111001101001001011011011	;
		random_num_table[28]  <= 32'b	00000100000100001110100011010100	;
		random_num_table[29]  <= 32'b	00011011010010100110111001011100	;
		random_num_table[30]  <= 32'b	00001111110111011010110011100001	;
		random_num_table[31]  <= 32'b	00001010011001100110101010100100	;
		random_num_table[32]  <= 32'b	00010111100101101011001011100100	;
		random_num_table[33]  <= 32'b	00001011100111011100100110100101	;
		random_num_table[34]  <= 32'b	00011101110011100111000111000110	;
		random_num_table[35]  <= 32'b	00010101101011110100101101011110	;
		random_num_table[36]  <= 32'b	00011110010001110100001010101001	;
		random_num_table[37]  <= 32'b	00000000001000110010101100101100	;
		random_num_table[38]  <= 32'b	00001111110000000010001111100001	;
		random_num_table[39]  <= 32'b	00010111001101010000110001010101	;
		random_num_table[40]  <= 32'b	00010100011001100111010001000101	;
		random_num_table[41]  <= 32'b	00011100111101001100110001001011	;
		random_num_table[42]  <= 32'b	00001011001110111010101100011000	;
		random_num_table[43]  <= 32'b	00001000110101010110011000000010	;
		random_num_table[44]  <= 32'b	00001000101101011000010111101101	;
		random_num_table[45]  <= 32'b	00010011011110001001110010010000	;
		random_num_table[46]  <= 32'b	00011010101001100100000110101010	;
		random_num_table[47]  <= 32'b	00010100111110011010110110101111	;
		random_num_table[48]  <= 32'b	00010100111110010100101000101101	;
		random_num_table[49]  <= 32'b	00011010011110111000010110010111	;
		random_num_table[50]  <= 32'b	00001111110000000011000100011111	;
		random_num_table[51]  <= 32'b	00010110001000100001011110010000	;
		random_num_table[52]  <= 32'b	00000000100001000000111101100111	;
		random_num_table[53]  <= 32'b	00000010011001100011111111001110	;
		random_num_table[54]  <= 32'b	00000100001110000110110000100000	;
		random_num_table[55]  <= 32'b	00000000001100100000011100100111	;
		random_num_table[56]  <= 32'b	00010000010110010110110010110111	;
		random_num_table[57]  <= 32'b	00010100000111101000000001000101	;
		random_num_table[58]  <= 32'b	00011110111101111010011000100001	;
		random_num_table[59]  <= 32'b	00000010110100111110100111001100	;
		random_num_table[60]  <= 32'b	00010101100100110001000111110110	;
		random_num_table[61]  <= 32'b	00001011001111001100101001101000	;
		random_num_table[62]  <= 32'b	00011010101011100100011100001010	;
		random_num_table[63]  <= 32'b	00011100011110001000001100101101	;
		random_num_table[64]  <= 32'b	00001010011000000100001100010011	;
		random_num_table[65]  <= 32'b	00000010001111111111101100001010	;
		random_num_table[66]  <= 32'b	00011111110001100011110101011001	;
		random_num_table[67]  <= 32'b	00010100110001100110101010000100	;
		random_num_table[68]  <= 32'b	00000111000100000101111111110110	;
		random_num_table[69]  <= 32'b	00010001010111111011001110001100	;
		random_num_table[70]  <= 32'b	00011101011100110100011011011110	;
		random_num_table[71]  <= 32'b	00010100110010000100000010010101	;
		random_num_table[72]  <= 32'b	00011011000000010100000010110001	;
		random_num_table[73]  <= 32'b	00010000101100001000100001101000	;
		random_num_table[74]  <= 32'b	00011100010001010110001111110010	;
		random_num_table[75]  <= 32'b	00001010101000101110111001000110	;
		random_num_table[76]  <= 32'b	00000010000110100001010011111101	;
		random_num_table[77]  <= 32'b	00001101001011001100110000101010	;
		random_num_table[78]  <= 32'b	00010000010000000100011010011101	;
		random_num_table[79]  <= 32'b	00011001101100000001110010011011	;
		random_num_table[80]  <= 32'b	00001000100111110011000100101110	;
		random_num_table[81]  <= 32'b	00011111101011010010010011000111	;
		random_num_table[82]  <= 32'b	00000111110100110110010010111000	;
		random_num_table[83]  <= 32'b	00011100100000100011010010101011	;
		random_num_table[84]  <= 32'b	00001110001101111110110100000000	;
		random_num_table[85]  <= 32'b	00011100000101101111010010100011	;
		random_num_table[86]  <= 32'b	00010001010000111101111100100011	;
		random_num_table[87]  <= 32'b	00000111000101010011110100111010	;
		random_num_table[88]  <= 32'b	00001101011111100010000000011101	;
		random_num_table[89]  <= 32'b	00011001111010110101010010111110	;
		random_num_table[90]  <= 32'b	00011010010010000101110011101010	;
		random_num_table[91]  <= 32'b	00001111101100000101100011101100	;
		random_num_table[92]  <= 32'b	00011111000011111110100111000101	;
		random_num_table[93]  <= 32'b	00001010001100111100101001111100	;
		random_num_table[94]  <= 32'b	00010011010100010100000011011100	;
		random_num_table[95]  <= 32'b	00011001010000001001101011100110	;
		random_num_table[96]  <= 32'b	00000010001001010010010001101100	;
		random_num_table[97]  <= 32'b	00001001001101100001111010100111	;
		random_num_table[98]  <= 32'b	00011001010010100011010001001100	;
		random_num_table[99]  <= 32'b	00011110011011001110000000001110	;
		random_num_table[100]  <= 32'b	00001000000110101110011101010010	;
		random_num_table[101]  <= 32'b	00001100001110010111011001100001	;
		random_num_table[102]  <= 32'b	00001010011100000001011101111001	;
		random_num_table[103]  <= 32'b	00000101100011010001111001111110	;
		random_num_table[104]  <= 32'b	00000010101100101011101101011000	;
		random_num_table[105]  <= 32'b	00011110000011101100101110110010	;
		random_num_table[106]  <= 32'b	00001100011011110001101010110111	;
		random_num_table[107]  <= 32'b	00000011110011111010100110110010	;
		random_num_table[108]  <= 32'b	00010100111101001110001110111100	;
		random_num_table[109]  <= 32'b	00000101001100111100100011001101	;
		random_num_table[110]  <= 32'b	00011101111101111110001100101110	;
		random_num_table[111]  <= 32'b	00001101111011111111111111101111	;
		random_num_table[112]  <= 32'b	00011011001001100101111101010101	;
		random_num_table[113]  <= 32'b	00010110011110011100011101001001	;
		random_num_table[114]  <= 32'b	00011010101101000010010000100000	;
		random_num_table[115]  <= 32'b	00000100100101011011111010110111	;
		random_num_table[116]  <= 32'b	00000010100001101010111100000010	;
		random_num_table[117]  <= 32'b	00001010010100011100110100010110	;
		random_num_table[118]  <= 32'b	00001101111000011010110100000001	;
		random_num_table[119]  <= 32'b	00000111011111101010011110111010	;
		random_num_table[120]  <= 32'b	00010100010100111010110011010001	;
		random_num_table[121]  <= 32'b	00011100000111001110111100001011	;
		random_num_table[122]  <= 32'b	00000011110110111100100100000100	;
		random_num_table[123]  <= 32'b	00001100010110011100111000110100	;
		random_num_table[124]  <= 32'b	00011101001111010110000100100010	;
		random_num_table[125]  <= 32'b	00000000001010000011101110100101	;
		random_num_table[126]  <= 32'b	00000010100010010100110110100000	;
		random_num_table[127]  <= 32'b	00000111110101111101000000001110	;
		random_num_table[128]  <= 32'b	00010001110001010001010000101110	;
		random_num_table[129]  <= 32'b	00000011001101101001101100100010	;
		random_num_table[130]  <= 32'b	00000110100100111110001011000011	;
		random_num_table[131]  <= 32'b	00001100000000001110001100100011	;
		random_num_table[132]  <= 32'b	00001000100100010101010000000010	;
		random_num_table[133]  <= 32'b	00000101000011100111101011111111	;
		random_num_table[134]  <= 32'b	00001011101010000100000100011101	;
		random_num_table[135]  <= 32'b	00001111010011101111101001010101	;
		random_num_table[136]  <= 32'b	00010101111110011111011101100101	;
		random_num_table[137]  <= 32'b	00010101001100000011101111100100	;
		random_num_table[138]  <= 32'b	00011110110000010000111101101011	;
		random_num_table[139]  <= 32'b	00010000010101100100001011110110	;
		random_num_table[140]  <= 32'b	00001110001010100101010110100110	;
		random_num_table[141]  <= 32'b	00010100100010010101000011010111	;
		random_num_table[142]  <= 32'b	00010111001100110111011110010001	;
		random_num_table[143]  <= 32'b	00000001000001000101010010110101	;
		random_num_table[144]  <= 32'b	00010011000000011101000001100110	;
		random_num_table[145]  <= 32'b	00010000100111110001111011010011	;
		random_num_table[146]  <= 32'b	00001110101011111111101000111110	;
		random_num_table[147]  <= 32'b	00010100101110100010001010000100	;
		random_num_table[148]  <= 32'b	00000111001101110111011011000000	;
		random_num_table[149]  <= 32'b	00011111000010011100010011110101	;
		random_num_table[150]  <= 32'b	00000011001111011101011111001010	;
		random_num_table[151]  <= 32'b	00011011111001100010001010010110	;
		random_num_table[152]  <= 32'b	00011100110100111011010011101110	;
		random_num_table[153]  <= 32'b	00000110111010011110111100000100	;
		random_num_table[154]  <= 32'b	00001101011101000011011001100011	;
		random_num_table[155]  <= 32'b	00010010000100101010111011011111	;
		random_num_table[156]  <= 32'b	00000011101011101010101111111100	;
		random_num_table[157]  <= 32'b	00000010001111001001111100100001	;
		random_num_table[158]  <= 32'b	00011001000011111000111110100111	;
		random_num_table[159]  <= 32'b	00011011010001010010101000001000	;
		random_num_table[160]  <= 32'b	00000001100010011111110011111011	;
		random_num_table[161]  <= 32'b	00001000010101000100010001110011	;
		random_num_table[162]  <= 32'b	00010001111110011110010101101110	;
		random_num_table[163]  <= 32'b	00010001111001100011001001011000	;
		random_num_table[164]  <= 32'b	00000110000010111000110001010000	;
		random_num_table[165]  <= 32'b	00011111010111001110110101100101	;
		random_num_table[166]  <= 32'b	00000010011100010101000101100110	;
		random_num_table[167]  <= 32'b	00011101000110111000011001000110	;
		random_num_table[168]  <= 32'b	00011000100010101010110100101011	;
		random_num_table[169]  <= 32'b	00011011101011111000000001000010	;
		random_num_table[170]  <= 32'b	00000000010000111010001000000011	;
		random_num_table[171]  <= 32'b	00010001011101010000000110010111	;
		random_num_table[172]  <= 32'b	00010100011000010110010010110010	;
		random_num_table[173]  <= 32'b	00001101101000110011001011000101	;
		random_num_table[174]  <= 32'b	00000011110101110010001100010100	;
		random_num_table[175]  <= 32'b	00011100101010110000100010101011	;
		random_num_table[176]  <= 32'b	00010001000011100101001011100111	;
		random_num_table[177]  <= 32'b	00000111101001010000111110101100	;
		random_num_table[178]  <= 32'b	00000010111110000111010100111011	;
		random_num_table[179]  <= 32'b	00010101111101101110100001110101	;
		random_num_table[180]  <= 32'b	00011111101111010101111010101110	;
		random_num_table[181]  <= 32'b	00000101111101111000100100010000	;
		random_num_table[182]  <= 32'b	00001011101101001110111000010000	;
		random_num_table[183]  <= 32'b	00011110001101011100001001101000	;
		random_num_table[184]  <= 32'b	00000101110011100010011000101001	;
		random_num_table[185]  <= 32'b	00000110100000010011001111011011	;
		random_num_table[186]  <= 32'b	00011100101000110111010110011101	;
		random_num_table[187]  <= 32'b	00011110101010110000100011001000	;
		random_num_table[188]  <= 32'b	00010101110011011111001110010001	;
		random_num_table[189]  <= 32'b	00000000010100011100010000100110	;
		random_num_table[190]  <= 32'b	00001111001010011000110011011111	;
		random_num_table[191]  <= 32'b	00010010111101000101110010001101	;
		random_num_table[192]  <= 32'b	00000011100001001010011000111001	;
		random_num_table[193]  <= 32'b	00000010000011011101100011000010	;
		random_num_table[194]  <= 32'b	00000111011000101101101110001001	;
		random_num_table[195]  <= 32'b	00011111100100001010110011000010	;
		random_num_table[196]  <= 32'b	00001000101001101111011000101100	;
		random_num_table[197]  <= 32'b	00001100110111110110101010001001	;
		random_num_table[198]  <= 32'b	00000010100010010111000110100010	;
		random_num_table[199]  <= 32'b	00000011000001010010010100100011	;
		random_num_table[200]  <= 32'b	00011100010100111110101001010110	;
		random_num_table[201]  <= 32'b	00000110101011101011001101111010	;
		random_num_table[202]  <= 32'b	00001000111101001110001100010000	;
		random_num_table[203]  <= 32'b	00011000011101101111000010101101	;
		random_num_table[204]  <= 32'b	00011110011100010000011001101100	;
		random_num_table[205]  <= 32'b	00010101100001110110000110110011	;
		random_num_table[206]  <= 32'b	00010110001100010000100110110010	;
		random_num_table[207]  <= 32'b	00000110100111101010101100110011	;
		random_num_table[208]  <= 32'b	00001000001101110101100001101000	;
		random_num_table[209]  <= 32'b	00001000000100010000000001110010	;
		random_num_table[210]  <= 32'b	00010001001110110111101100011100	;
		random_num_table[211]  <= 32'b	00010010111000001111101100001000	;
		random_num_table[212]  <= 32'b	00011001101011101101000011100110	;
		random_num_table[213]  <= 32'b	00011011101000000100001001110101	;
		random_num_table[214]  <= 32'b	00001100100100110110101001111110	;
		random_num_table[215]  <= 32'b	00001101111100100000101000011001	;
		random_num_table[216]  <= 32'b	00001000110111111100011011001101	;
		random_num_table[217]  <= 32'b	00001110110110110111110110001010	;
		random_num_table[218]  <= 32'b	00011100000110111011110000100111	;
		random_num_table[219]  <= 32'b	00010001010100000000100010101001	;
		random_num_table[220]  <= 32'b	00001101100101101001101101000110	;
		random_num_table[221]  <= 32'b	00011100100110011011011101001000	;
		random_num_table[222]  <= 32'b	00000011000010011111000000000010	;
		random_num_table[223]  <= 32'b	00010110100011000000111111011010	;
		random_num_table[224]  <= 32'b	00000111100001011101110100001011	;
		random_num_table[225]  <= 32'b	00001001111011100100110010011101	;
		random_num_table[226]  <= 32'b	00000100010010111001001010100000	;
		random_num_table[227]  <= 32'b	00000011111010000100101001000110	;
		random_num_table[228]  <= 32'b	00001110101001111001110111110010	;
		random_num_table[229]  <= 32'b	00000010011010110101100101111011	;
		random_num_table[230]  <= 32'b	00011101000100101000010000100101	;
		random_num_table[231]  <= 32'b	00010001100011001000101010000011	;
		random_num_table[232]  <= 32'b	00001011111010001000011111111000	;
		random_num_table[233]  <= 32'b	00000100101001110111001000000110	;
		random_num_table[234]  <= 32'b	00000010011110100000011111001001	;
		random_num_table[235]  <= 32'b	00000100100110100000011010100011	;
		random_num_table[236]  <= 32'b	00011100110001000111101000001111	;
		random_num_table[237]  <= 32'b	00011111000100011110010001001000	;
		random_num_table[238]  <= 32'b	00001100100001110101101110101110	;
		random_num_table[239]  <= 32'b	00010001110000111111000101101101	;
		random_num_table[240]  <= 32'b	00001001100111110001000110110100	;
		random_num_table[241]  <= 32'b	00000000010101110000111111111010	;
		random_num_table[242]  <= 32'b	00010011000100100101111101101111	;
		random_num_table[243]  <= 32'b	00000111111111101001110011000000	;
		random_num_table[244]  <= 32'b	00000110101010111101110000001011	;
		random_num_table[245]  <= 32'b	00001010001011100111111110000110	;
		random_num_table[246]  <= 32'b	00000101100010110011111010000110	;
		random_num_table[247]  <= 32'b	00010101100001011101011000010100	;
		random_num_table[248]  <= 32'b	00011010110011011110001010100001	;
		random_num_table[249]  <= 32'b	00001010000111100010010000001111	;
		random_num_table[250]  <= 32'b	00011010101101010110111100001100	;
		random_num_table[251]  <= 32'b	00011011110010010111010010010110	;
		random_num_table[252]  <= 32'b	00011011111001100110010011011100	;
		random_num_table[253]  <= 32'b	00010101001111011001000000001011	;
		random_num_table[254]  <= 32'b	00010010110111011111110100010111	;
		random_num_table[255]  <= 32'b	00001000000001110011011000110010	;			
	end
endmodule
