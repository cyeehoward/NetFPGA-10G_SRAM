`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:43:16 01/19/2015 
// Design Name: 
// Module Name:    rand_table_1 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module rand_table_1(axi_aclk , axi_aresetn , index_num , rand_out , en);
	input			axi_aclk , axi_aresetn , en;
	input		[7:0]	index_num;
	output		[31:0]	rand_out;

	reg 		[31:0]	random_num_table  [255:0];

	assign rand_out = en?random_num_table[index_num]:32'd0;
	
	always@(posedge axi_aclk)
	begin
		random_num_table[0]  <= 32'b	00011111011001010111011011010011	;
		random_num_table[1]  <= 32'b	00011110001010111110111100101101	;
		random_num_table[2]  <= 32'b	00000001110001111001001001100011	;
		random_num_table[3]  <= 32'b	00000010000110111001101101110101	;
		random_num_table[4]  <= 32'b	00000000010011011101111000111011	;
		random_num_table[5]  <= 32'b	00010111000101011101001010010101	;
		random_num_table[6]  <= 32'b	00010100111011001101100011001010	;
		random_num_table[7]  <= 32'b	00010101001011001101001101101100	;
		random_num_table[8]  <= 32'b	00010101010100000001010011011011	;
		random_num_table[9]  <= 32'b	00010000001111001011010101011100	;
		random_num_table[10]  <= 32'b	00010010111011101110111111011110	;
		random_num_table[11]  <= 32'b	00011000111011111010101010100001	;
		random_num_table[12]  <= 32'b	00001101100011001111100100001110	;
		random_num_table[13]  <= 32'b	00000011000011000110100001101111	;
		random_num_table[14]  <= 32'b	00010011100010100100001110101100	;
		random_num_table[15]  <= 32'b	00000101001111000011011001011011	;
		random_num_table[16]  <= 32'b	00011010001000010011010010101110	;
		random_num_table[17]  <= 32'b	00000111111011000111000010110010	;
		random_num_table[18]  <= 32'b	00011010010100101101110110001011	;
		random_num_table[19]  <= 32'b	00000010111100101100111111110001	;
		random_num_table[20]  <= 32'b	00001011010101010000110101011100	;
		random_num_table[21]  <= 32'b	00001011111111101001000100001111	;
		random_num_table[22]  <= 32'b	00000011011100011100001101001100	;
		random_num_table[23]  <= 32'b	00001011110110011111000011110011	;
		random_num_table[24]  <= 32'b	00001101000011011110111001110010	;
		random_num_table[25]  <= 32'b	00000111000111010010011010111000	;
		random_num_table[26]  <= 32'b	00000010100001110111001101101010	;
		random_num_table[27]  <= 32'b	00001001010001111011011100000011	;
		random_num_table[28]  <= 32'b	00011100100000110000011000010000	;
		random_num_table[29]  <= 32'b	00001011010110101001010110000110	;
		random_num_table[30]  <= 32'b	00001011100010101111000011101110	;
		random_num_table[31]  <= 32'b	00000101110011010000111111111100	;
		random_num_table[32]  <= 32'b	00001101001000110000100011101111	;
		random_num_table[33]  <= 32'b	00010011100001110011101000000000	;
		random_num_table[34]  <= 32'b	00000011111010110011101101011001	;
		random_num_table[35]  <= 32'b	00001101000001011011011000001000	;
		random_num_table[36]  <= 32'b	00000101110101010101011100000001	;
		random_num_table[37]  <= 32'b	00010010101010000010110110100100	;
		random_num_table[38]  <= 32'b	00011111010110000010101101100010	;
		random_num_table[39]  <= 32'b	00000110101110101001111011010011	;
		random_num_table[40]  <= 32'b	00001010110001001001011110100001	;
		random_num_table[41]  <= 32'b	00010101100111101011100011011000	;
		random_num_table[42]  <= 32'b	00010011010111100101011111111001	;
		random_num_table[43]  <= 32'b	00011100001100001100111110011110	;
		random_num_table[44]  <= 32'b	00001101110001111100001101111101	;
		random_num_table[45]  <= 32'b	00011110001000010011111101110001	;
		random_num_table[46]  <= 32'b	00010111101101010110011001111001	;
		random_num_table[47]  <= 32'b	00000111000011010001000011001001	;
		random_num_table[48]  <= 32'b	00001101010101111000111100000000	;
		random_num_table[49]  <= 32'b	00011011110111011010000000000101	;
		random_num_table[50]  <= 32'b	00000111101011000100101100010011	;
		random_num_table[51]  <= 32'b	00000001110101000010100000001110	;
		random_num_table[52]  <= 32'b	00010011011010110110010011110110	;
		random_num_table[53]  <= 32'b	00011001100000011011000110011100	;
		random_num_table[54]  <= 32'b	00000111011100101111110000110001	;
		random_num_table[55]  <= 32'b	00011011100010001111010111101111	;
		random_num_table[56]  <= 32'b	00010010010100100001100110011101	;
		random_num_table[57]  <= 32'b	00001101100001011110010111110010	;
		random_num_table[58]  <= 32'b	00000001011100000011011011100010	;
		random_num_table[59]  <= 32'b	00001110000111011100011110101001	;
		random_num_table[60]  <= 32'b	00011010100100101111111000101010	;
		random_num_table[61]  <= 32'b	00011111000001111010001100011111	;
		random_num_table[62]  <= 32'b	00000011010101000100100100001011	;
		random_num_table[63]  <= 32'b	00011100000001010100101110101111	;
		random_num_table[64]  <= 32'b	00001100101101111010000011111011	;
		random_num_table[65]  <= 32'b	00000001011010011010000000111110	;
		random_num_table[66]  <= 32'b	00010100111100111000010000001001	;
		random_num_table[67]  <= 32'b	00000001000110100110111111010111	;
		random_num_table[68]  <= 32'b	00010011111010111001000011110101	;
		random_num_table[69]  <= 32'b	00000101010110011010011100101011	;
		random_num_table[70]  <= 32'b	00001001011111010010011101001001	;
		random_num_table[71]  <= 32'b	00010011110001011111101011100010	;
		random_num_table[72]  <= 32'b	00010001011000100100100010101111	;
		random_num_table[73]  <= 32'b	00001110010101101010001010010001	;
		random_num_table[74]  <= 32'b	00010000000101000100001001010011	;
		random_num_table[75]  <= 32'b	00000001111011110110010001110110	;
		random_num_table[76]  <= 32'b	00010001101110001110001011001000	;
		random_num_table[77]  <= 32'b	00011110001110111101111000010000	;
		random_num_table[78]  <= 32'b	00010111000110100110011001100100	;
		random_num_table[79]  <= 32'b	00000000111001110111101110101010	;
		random_num_table[80]  <= 32'b	00001001011111011011001000000001	;
		random_num_table[81]  <= 32'b	00011110001100111100011100111000	;
		random_num_table[82]  <= 32'b	00010111011101111111100111100101	;
		random_num_table[83]  <= 32'b	00010000101000110111011000101101	;
		random_num_table[84]  <= 32'b	00010011101101000001101001111011	;
		random_num_table[85]  <= 32'b	00011010010100101011000000000110	;
		random_num_table[86]  <= 32'b	00000110110101001110001100110100	;
		random_num_table[87]  <= 32'b	00011100011100011000000100000011	;
		random_num_table[88]  <= 32'b	00010010101110001001101111110110	;
		random_num_table[89]  <= 32'b	00010100011101011011100001011001	;
		random_num_table[90]  <= 32'b	00000011010011010001000110010101	;
		random_num_table[91]  <= 32'b	00000101001001001100001000110001	;
		random_num_table[92]  <= 32'b	00000010001010010000101001100111	;
		random_num_table[93]  <= 32'b	00001000101011001010100111010110	;
		random_num_table[94]  <= 32'b	00001100100001000011101000110110	;
		random_num_table[95]  <= 32'b	00001111110010111111000011010010	;
		random_num_table[96]  <= 32'b	00011101110100010010100000000001	;
		random_num_table[97]  <= 32'b	00010001100011000000111011110110	;
		random_num_table[98]  <= 32'b	00011011101110100101001011011010	;
		random_num_table[99]  <= 32'b	00010101100111111000100111101100	;
		random_num_table[100]  <= 32'b	00001001100101101111100001001110	;
		random_num_table[101]  <= 32'b	00011000000110110001010110000100	;
		random_num_table[102]  <= 32'b	00010010011100000101101010011001	;
		random_num_table[103]  <= 32'b	00000111010000011101011011101100	;
		random_num_table[104]  <= 32'b	00011011101011000001011111110001	;
		random_num_table[105]  <= 32'b	00011101001101011101011000101110	;
		random_num_table[106]  <= 32'b	00010111101011110110111111101101	;
		random_num_table[107]  <= 32'b	00011100111110010101011110001001	;
		random_num_table[108]  <= 32'b	00001100001001111000010010110010	;
		random_num_table[109]  <= 32'b	00001010100100000000110000010011	;
		random_num_table[110]  <= 32'b	00001101100110111110100100111111	;
		random_num_table[111]  <= 32'b	00001011111111000111001010101111	;
		random_num_table[112]  <= 32'b	00001101110100101101101000001101	;
		random_num_table[113]  <= 32'b	00011000111001100011000110011011	;
		random_num_table[114]  <= 32'b	00001100101110010100111110101001	;
		random_num_table[115]  <= 32'b	00001001010111110110001010101001	;
		random_num_table[116]  <= 32'b	00001010101001110111101000000001	;
		random_num_table[117]  <= 32'b	00010001100011000010001000100011	;
		random_num_table[118]  <= 32'b	00010000010010101010111000010101	;
		random_num_table[119]  <= 32'b	00001100001111110100110011111101	;
		random_num_table[120]  <= 32'b	00000001010011100000001101110000	;
		random_num_table[121]  <= 32'b	00000110011111011000010100111101	;
		random_num_table[122]  <= 32'b	00000110110110110100010100100001	;
		random_num_table[123]  <= 32'b	00000100000011000100101100110111	;
		random_num_table[124]  <= 32'b	00010010100000000110111000000001	;
		random_num_table[125]  <= 32'b	00000110110010111000110000101111	;
		random_num_table[126]  <= 32'b	00010010001101010010001101111101	;
		random_num_table[127]  <= 32'b	00011110101000010100110111001000	;
		random_num_table[128]  <= 32'b	00001011110000101000110101010000	;
		random_num_table[129]  <= 32'b	00010110001011011111010111010001	;
		random_num_table[130]  <= 32'b	00011110011101100010010111011000	;
		random_num_table[131]  <= 32'b	00011011011011010100100100011010	;
		random_num_table[132]  <= 32'b	00001010100110101101100101000111	;
		random_num_table[133]  <= 32'b	00001000010111010101000100000111	;
		random_num_table[134]  <= 32'b	00011011000011110101000000111001	;
		random_num_table[135]  <= 32'b	00001100011001011001010110000010	;
		random_num_table[136]  <= 32'b	00010011100100000100000010100111	;
		random_num_table[137]  <= 32'b	00001101010100001101110101011110	;
		random_num_table[138]  <= 32'b	00001010100000101101010111000010	;
		random_num_table[139]  <= 32'b	00011010000011111110011100100100	;
		random_num_table[140]  <= 32'b	00001101001000110110111111100010	;
		random_num_table[141]  <= 32'b	00011111000101011010100011000111	;
		random_num_table[142]  <= 32'b	00001011100011100010010101111010	;
		random_num_table[143]  <= 32'b	00010100000111101101100100101100	;
		random_num_table[144]  <= 32'b	00011000101110001011111110011111	;
		random_num_table[145]  <= 32'b	00011100000111100101001000011101	;
		random_num_table[146]  <= 32'b	00000100101111100111011101011101	;
		random_num_table[147]  <= 32'b	00010011101110000000100000110000	;
		random_num_table[148]  <= 32'b	00000101000011100010001010000000	;
		random_num_table[149]  <= 32'b	00000000101000001011000110100110	;
		random_num_table[150]  <= 32'b	00001011100110110000010010011111	;
		random_num_table[151]  <= 32'b	00000001001111101100000111010111	;
		random_num_table[152]  <= 32'b	00001001100001001110010111011101	;
		random_num_table[153]  <= 32'b	00000101110111011101101111100010	;
		random_num_table[154]  <= 32'b	00000110001001101000010111111110	;
		random_num_table[155]  <= 32'b	00010100111101111110001111101010	;
		random_num_table[156]  <= 32'b	00001101010000001000101000110011	;
		random_num_table[157]  <= 32'b	00000010011101000111010100001100	;
		random_num_table[158]  <= 32'b	00000001000111010100111010011010	;
		random_num_table[159]  <= 32'b	00001111001101111000011110111111	;
		random_num_table[160]  <= 32'b	00000000011010010111111101110101	;
		random_num_table[161]  <= 32'b	00001100010100111111100100010100	;
		random_num_table[162]  <= 32'b	00010101110100011100011001010111	;
		random_num_table[163]  <= 32'b	00010011110001010001000100010101	;
		random_num_table[164]  <= 32'b	00011010001100011011101111110101	;
		random_num_table[165]  <= 32'b	00000101110111000000111100001000	;
		random_num_table[166]  <= 32'b	00011111110000001101100111101000	;
		random_num_table[167]  <= 32'b	00011011011001001001111100010000	;
		random_num_table[168]  <= 32'b	00000001010100110110010010101001	;
		random_num_table[169]  <= 32'b	00011110100100101111110101011110	;
		random_num_table[170]  <= 32'b	00011110010000011100000001001101	;
		random_num_table[171]  <= 32'b	00001111111111000100110011111001	;
		random_num_table[172]  <= 32'b	00000010110000101101011010010100	;
		random_num_table[173]  <= 32'b	00000011110011011111011000011010	;
		random_num_table[174]  <= 32'b	00010001001011110101010001100011	;
		random_num_table[175]  <= 32'b	00011101011100001001010100101010	;
		random_num_table[176]  <= 32'b	00001110111101110010010011111001	;
		random_num_table[177]  <= 32'b	00000101011110100010011101101111	;
		random_num_table[178]  <= 32'b	00011000111000011000101000101001	;
		random_num_table[179]  <= 32'b	00010110100100001110101001100101	;
		random_num_table[180]  <= 32'b	00001001110010101010011011001100	;
		random_num_table[181]  <= 32'b	00001101100101011101000011101110	;
		random_num_table[182]  <= 32'b	00001010100011111111110010111111	;
		random_num_table[183]  <= 32'b	00001101101000010110010011110010	;
		random_num_table[184]  <= 32'b	00011111101111100001010100100011	;
		random_num_table[185]  <= 32'b	00010010101110011110110001101101	;
		random_num_table[186]  <= 32'b	00001101101011111001111110011001	;
		random_num_table[187]  <= 32'b	00011010110010000001110000100100	;
		random_num_table[188]  <= 32'b	00010011111101011001101001101110	;
		random_num_table[189]  <= 32'b	00010101011000111111100001000110	;
		random_num_table[190]  <= 32'b	00000110000110010010001000111011	;
		random_num_table[191]  <= 32'b	00000110010100100111110011110001	;
		random_num_table[192]  <= 32'b	00011011110100001100011001000010	;
		random_num_table[193]  <= 32'b	00000011100110010010001011101110	;
		random_num_table[194]  <= 32'b	00010001001101000011100011011001	;
		random_num_table[195]  <= 32'b	00011001100110110101001010110000	;
		random_num_table[196]  <= 32'b	00010011010010111011010010000111	;
		random_num_table[197]  <= 32'b	00010010000000010001010110000010	;
		random_num_table[198]  <= 32'b	00010100010010001110001010000010	;
		random_num_table[199]  <= 32'b	00000011111011110110110000001001	;
		random_num_table[200]  <= 32'b	00001011000111011010111101110010	;
		random_num_table[201]  <= 32'b	00011000100010111001010001001001	;
		random_num_table[202]  <= 32'b	00001100011111100100111111000011	;
		random_num_table[203]  <= 32'b	00001001000011000100000101101010	;
		random_num_table[204]  <= 32'b	00001010001110011010101011011110	;
		random_num_table[205]  <= 32'b	00011111101010010001011100111011	;
		random_num_table[206]  <= 32'b	00011001111101001100100101011010	;
		random_num_table[207]  <= 32'b	00000001011011111001101001010101	;
		random_num_table[208]  <= 32'b	00010111111101100100001100101111	;
		random_num_table[209]  <= 32'b	00010101100010010000110011110010	;
		random_num_table[210]  <= 32'b	00001001010010011011110111011001	;
		random_num_table[211]  <= 32'b	00010001111010001010100010001100	;
		random_num_table[212]  <= 32'b	00001111100010010100100100111000	;
		random_num_table[213]  <= 32'b	00001110101110010011010001011101	;
		random_num_table[214]  <= 32'b	00010001000111100010101110111101	;
		random_num_table[215]  <= 32'b	00001000101110011111101111101000	;
		random_num_table[216]  <= 32'b	00001001100000001010001100010100	;
		random_num_table[217]  <= 32'b	00011001111001010111001011100111	;
		random_num_table[218]  <= 32'b	00001001110001110111000101111000	;
		random_num_table[219]  <= 32'b	00000100011101000000101011001100	;
		random_num_table[220]  <= 32'b	00000111100010110101101011111110	;
		random_num_table[221]  <= 32'b	00000010111111100011011011000101	;
		random_num_table[222]  <= 32'b	00000001001110001111001100101011	;
		random_num_table[223]  <= 32'b	00010110000010110100111001010010	;
		random_num_table[224]  <= 32'b	00011100011100111100001100000010	;
		random_num_table[225]  <= 32'b	00010110110001011010001011101011	;
		random_num_table[226]  <= 32'b	00011111100001110000011110000110	;
		random_num_table[227]  <= 32'b	00011100011110100110010100001111	;
		random_num_table[228]  <= 32'b	00011000010101110010000110101010	;
		random_num_table[229]  <= 32'b	00010010111001001000100011011010	;
		random_num_table[230]  <= 32'b	00010000100001001001011110001011	;
		random_num_table[231]  <= 32'b	00011101000100011110100111101100	;
		random_num_table[232]  <= 32'b	00010000001000011001001011101111	;
		random_num_table[233]  <= 32'b	00011000100101000101100011011100	;
		random_num_table[234]  <= 32'b	00001100000111110010110101110000	;
		random_num_table[235]  <= 32'b	00000011000111110100001001101001	;
		random_num_table[236]  <= 32'b	00000111010111010011111000011010	;
		random_num_table[237]  <= 32'b	00001110010001001100001011000110	;
		random_num_table[238]  <= 32'b	00010111111011011011111111111001	;
		random_num_table[239]  <= 32'b	00011000100111011101101010011101	;
		random_num_table[240]  <= 32'b	00010110011011001100110001010100	;
		random_num_table[241]  <= 32'b	00000000101100011111010111110100	;
		random_num_table[242]  <= 32'b	00010111101110110010100110010110	;
		random_num_table[243]  <= 32'b	00000100111001001110111111011101	;
		random_num_table[244]  <= 32'b	00011001001100100101001011011100	;
		random_num_table[245]  <= 32'b	00010000100110100101010010110101	;
		random_num_table[246]  <= 32'b	00011111010001011111101000000100	;
		random_num_table[247]  <= 32'b	00001110000101111111100010000010	;
		random_num_table[248]  <= 32'b	00011010100110010101001011100000	;
		random_num_table[249]  <= 32'b	00001101111011100000001010111111	;
		random_num_table[250]  <= 32'b	00011010101110000100100100110010	;
		random_num_table[251]  <= 32'b	00001101100110001101101100100100	;
		random_num_table[252]  <= 32'b	00001010000000110100110000001100	;
		random_num_table[253]  <= 32'b	00001101010111100111001101110010	;
		random_num_table[254]  <= 32'b	00001111111101101001011110100100	;
		random_num_table[255]  <= 32'b	00010000110000011101101010001100	;
	end
endmodule
