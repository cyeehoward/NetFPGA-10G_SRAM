`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:54:32 01/19/2015 
// Design Name: 
// Module Name:    rand_table_5 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module rand_table_5(axi_aclk , axi_aresetn , index_num , rand_out , en);
	input			axi_aclk , axi_aresetn , en;
	input		[7:0]	index_num;
	output		[31:0]	rand_out;

	reg 		[31:0]	random_num_table  [255:0];

	assign rand_out = en?random_num_table[index_num]:32'd0;
	
	always@(posedge axi_aclk)
	begin
		random_num_table[0]  <= 32'b	00010101011110110001111000110011	;
		random_num_table[1]  <= 32'b	00000101100100110011011100011011	;
		random_num_table[2]  <= 32'b	00000100000010101000001010001011	;
		random_num_table[3]  <= 32'b	00010111111000011011000000011000	;
		random_num_table[4]  <= 32'b	00010010101100011001110100110110	;
		random_num_table[5]  <= 32'b	00000111111110000111101110001010	;
		random_num_table[6]  <= 32'b	00011101111010011001010010110111	;
		random_num_table[7]  <= 32'b	00011011101100010100110000011000	;
		random_num_table[8]  <= 32'b	00011101100111101010000001011001	;
		random_num_table[9]  <= 32'b	00010111001110010000110011011001	;
		random_num_table[10]  <= 32'b	00001000100101001011011110001101	;
		random_num_table[11]  <= 32'b	00011111111110100011011100111101	;
		random_num_table[12]  <= 32'b	00010101000011011111110111010011	;
		random_num_table[13]  <= 32'b	00010100011011000111000100111001	;
		random_num_table[14]  <= 32'b	00010001111101011011010001010111	;
		random_num_table[15]  <= 32'b	00011001111000011010011011110100	;
		random_num_table[16]  <= 32'b	00000000101000101000101101001000	;
		random_num_table[17]  <= 32'b	00010100011001101000100110100011	;
		random_num_table[18]  <= 32'b	00001001001001010000001001110100	;
		random_num_table[19]  <= 32'b	00011000110110000001100101110101	;
		random_num_table[20]  <= 32'b	00011110010111000000111101110010	;
		random_num_table[21]  <= 32'b	00010101100001010010101100010011	;
		random_num_table[22]  <= 32'b	00000000100000100010101100111010	;
		random_num_table[23]  <= 32'b	00010111010100101010001000101110	;
		random_num_table[24]  <= 32'b	00000011000011010010110110110010	;
		random_num_table[25]  <= 32'b	00001011011011011110101011011111	;
		random_num_table[26]  <= 32'b	00001110001110001101110110111010	;
		random_num_table[27]  <= 32'b	00011010001001101111100101100100	;
		random_num_table[28]  <= 32'b	00001011111000010101011110100111	;
		random_num_table[29]  <= 32'b	00011000000000100000100110011000	;
		random_num_table[30]  <= 32'b	00001010010010000100101101001101	;
		random_num_table[31]  <= 32'b	00001100110100001100000011001100	;
		random_num_table[32]  <= 32'b	00000001101011001101000101001100	;
		random_num_table[33]  <= 32'b	00011110011010011110101101111011	;
		random_num_table[34]  <= 32'b	00001010100100001100111110111001	;
		random_num_table[35]  <= 32'b	00010100000011000101001010111011	;
		random_num_table[36]  <= 32'b	00011010011001001010011101110011	;
		random_num_table[37]  <= 32'b	00000100000111110010100001100011	;
		random_num_table[38]  <= 32'b	00001001101111100111000000101010	;
		random_num_table[39]  <= 32'b	00011011101001011111000101110110	;
		random_num_table[40]  <= 32'b	00000111010100010011000001010101	;
		random_num_table[41]  <= 32'b	00011001011100110000001100001001	;
		random_num_table[42]  <= 32'b	00000111000100101011001110111100	;
		random_num_table[43]  <= 32'b	00001011110000101101111000110111	;
		random_num_table[44]  <= 32'b	00011011100110100101101100010011	;
		random_num_table[45]  <= 32'b	00010111010100101101011101110100	;
		random_num_table[46]  <= 32'b	00000011001010011100111011111110	;
		random_num_table[47]  <= 32'b	00011011100011010111111000010001	;
		random_num_table[48]  <= 32'b	00001010011101001000110101011101	;
		random_num_table[49]  <= 32'b	00011101101110000110111010011001	;
		random_num_table[50]  <= 32'b	00001111110101001110011110101101	;
		random_num_table[51]  <= 32'b	00000110000110000111000000011010	;
		random_num_table[52]  <= 32'b	00001010100000100110010000010100	;
		random_num_table[53]  <= 32'b	00011000100101110100011000011100	;
		random_num_table[54]  <= 32'b	00000001110000011010110110000011	;
		random_num_table[55]  <= 32'b	00001100111000000100111000100001	;
		random_num_table[56]  <= 32'b	00001111001110110011010100011001	;
		random_num_table[57]  <= 32'b	00001010010011010010000110111010	;
		random_num_table[58]  <= 32'b	00001111011000101011001111001111	;
		random_num_table[59]  <= 32'b	00001010101110110100001101101100	;
		random_num_table[60]  <= 32'b	00011110111100111010011000110000	;
		random_num_table[61]  <= 32'b	00000100011111101011111100101010	;
		random_num_table[62]  <= 32'b	00010111110000100101110011110111	;
		random_num_table[63]  <= 32'b	00011001010010010100100010110111	;
		random_num_table[64]  <= 32'b	00001111001010101011010110011101	;
		random_num_table[65]  <= 32'b	00001100011101101101110001011110	;
		random_num_table[66]  <= 32'b	00001100101011111010011110001010	;
		random_num_table[67]  <= 32'b	00001010000010110001100011001010	;
		random_num_table[68]  <= 32'b	00000100100111100001000000111001	;
		random_num_table[69]  <= 32'b	00011000111010110110110101001010	;
		random_num_table[70]  <= 32'b	00000100100000011001001010010111	;
		random_num_table[71]  <= 32'b	00011101001110010101101011111011	;
		random_num_table[72]  <= 32'b	00010111010011101110110111110011	;
		random_num_table[73]  <= 32'b	00011101110110011100000011100100	;
		random_num_table[74]  <= 32'b	00000011001110011100010101000001	;
		random_num_table[75]  <= 32'b	00000010100101000000101000001011	;
		random_num_table[76]  <= 32'b	00011101010110001111111100010011	;
		random_num_table[77]  <= 32'b	00001001110100011111000010011001	;
		random_num_table[78]  <= 32'b	00001011001010100101001010100000	;
		random_num_table[79]  <= 32'b	00001010111011010011000110010111	;
		random_num_table[80]  <= 32'b	00001000001001110111010110000110	;
		random_num_table[81]  <= 32'b	00011011000111011010110001000011	;
		random_num_table[82]  <= 32'b	00010000001000110001000010010011	;
		random_num_table[83]  <= 32'b	00001010110110010101010110100111	;
		random_num_table[84]  <= 32'b	00000010100011001111001100000100	;
		random_num_table[85]  <= 32'b	00001111101111011111000101101101	;
		random_num_table[86]  <= 32'b	00010000010001010000110101000111	;
		random_num_table[87]  <= 32'b	00000000101110011010001000001001	;
		random_num_table[88]  <= 32'b	00001110001011001011100111000101	;
		random_num_table[89]  <= 32'b	00010010100100100110011111111110	;
		random_num_table[90]  <= 32'b	00010010100000011100100001101001	;
		random_num_table[91]  <= 32'b	00010111101111000111100111100111	;
		random_num_table[92]  <= 32'b	00000000011100111110010101000001	;
		random_num_table[93]  <= 32'b	00001010100100010000101101011111	;
		random_num_table[94]  <= 32'b	00000001111000011000110011111001	;
		random_num_table[95]  <= 32'b	00011001001001011010011111101000	;
		random_num_table[96]  <= 32'b	00001010111001010111000010010100	;
		random_num_table[97]  <= 32'b	00000010101001110101111101110011	;
		random_num_table[98]  <= 32'b	00011011100010011111001111100001	;
		random_num_table[99]  <= 32'b	00010101101110101011101101101011	;
		random_num_table[100]  <= 32'b	00011101111011110011100000011010	;
		random_num_table[101]  <= 32'b	00001000010101000111001110100100	;
		random_num_table[102]  <= 32'b	00010110110110011011010000110011	;
		random_num_table[103]  <= 32'b	00010011111011110010111010110101	;
		random_num_table[104]  <= 32'b	00001100001011110101101001001110	;
		random_num_table[105]  <= 32'b	00011100000111000110101010010000	;
		random_num_table[106]  <= 32'b	00000011011110010001001010001101	;
		random_num_table[107]  <= 32'b	00001000100110011000001101011010	;
		random_num_table[108]  <= 32'b	00000001110111111101101100001010	;
		random_num_table[109]  <= 32'b	00001011100011100101100100101010	;
		random_num_table[110]  <= 32'b	00011101011101001010111010011011	;
		random_num_table[111]  <= 32'b	00011011101101010111110010011101	;
		random_num_table[112]  <= 32'b	00001110010011011000011111101110	;
		random_num_table[113]  <= 32'b	00000111101101110100111111001100	;
		random_num_table[114]  <= 32'b	00011110100010111101010111011010	;
		random_num_table[115]  <= 32'b	00010101110010111111111111111001	;
		random_num_table[116]  <= 32'b	00000000101010010011101100010011	;
		random_num_table[117]  <= 32'b	00001001100110011111100110100111	;
		random_num_table[118]  <= 32'b	00001100000011011110110101100010	;
		random_num_table[119]  <= 32'b	00011001010010100101110001110000	;
		random_num_table[120]  <= 32'b	00011110011000010111111000010110	;
		random_num_table[121]  <= 32'b	00010101000000001010111001000001	;
		random_num_table[122]  <= 32'b	00011011001010101100100101000111	;
		random_num_table[123]  <= 32'b	00000011110001010011101010101000	;
		random_num_table[124]  <= 32'b	00000010000010010001110011001100	;
		random_num_table[125]  <= 32'b	00010101100101000011100111001010	;
		random_num_table[126]  <= 32'b	00001111000010111010001111100010	;
		random_num_table[127]  <= 32'b	00010011111011111010010010000000	;
		random_num_table[128]  <= 32'b	00011101111010000010000010010101	;
		random_num_table[129]  <= 32'b	00001100111110000100111111001000	;
		random_num_table[130]  <= 32'b	00011100011011000000001011100110	;
		random_num_table[131]  <= 32'b	00001110010101000001111000110000	;
		random_num_table[132]  <= 32'b	00010010100101101111010100000011	;
		random_num_table[133]  <= 32'b	00001110001010000011111001000100	;
		random_num_table[134]  <= 32'b	00000111001101111000010100011101	;
		random_num_table[135]  <= 32'b	00000111000101010001001110010010	;
		random_num_table[136]  <= 32'b	00011101110011101010101010010010	;
		random_num_table[137]  <= 32'b	00000000001110010100101101011100	;
		random_num_table[138]  <= 32'b	00000011000110110001010101001001	;
		random_num_table[139]  <= 32'b	00011111001010100110001001111100	;
		random_num_table[140]  <= 32'b	00000100111111010000110100110111	;
		random_num_table[141]  <= 32'b	00010111100101110001110101000010	;
		random_num_table[142]  <= 32'b	00011000111110111111010101001010	;
		random_num_table[143]  <= 32'b	00000001100101001110100111101010	;
		random_num_table[144]  <= 32'b	00001011010000111100011110101001	;
		random_num_table[145]  <= 32'b	00010101100001101010110100110000	;
		random_num_table[146]  <= 32'b	00011001001011011010010110110101	;
		random_num_table[147]  <= 32'b	00000101110110000001011001010011	;
		random_num_table[148]  <= 32'b	00010010101000011011100101011000	;
		random_num_table[149]  <= 32'b	00001011000100110110111100101010	;
		random_num_table[150]  <= 32'b	00001111101101110111100100100101	;
		random_num_table[151]  <= 32'b	00010101100011111111000010010110	;
		random_num_table[152]  <= 32'b	00001110010100111010011110100111	;
		random_num_table[153]  <= 32'b	00001101000101001101011011111001	;
		random_num_table[154]  <= 32'b	00000000011101100111101001111100	;
		random_num_table[155]  <= 32'b	00010011100001100111111011011000	;
		random_num_table[156]  <= 32'b	00001010010011110110001011101000	;
		random_num_table[157]  <= 32'b	00000111100010101100100001000111	;
		random_num_table[158]  <= 32'b	00011111101101101101000000100000	;
		random_num_table[159]  <= 32'b	00001010000011110110100110000010	;
		random_num_table[160]  <= 32'b	00010101100100111011010110011110	;
		random_num_table[161]  <= 32'b	00011110111111100100100100010110	;
		random_num_table[162]  <= 32'b	00001000001010010110010011110000	;
		random_num_table[163]  <= 32'b	00010101100001110110111111100110	;
		random_num_table[164]  <= 32'b	00011011000101011101110110000100	;
		random_num_table[165]  <= 32'b	00000110111111000111110001000001	;
		random_num_table[166]  <= 32'b	00010010101111010111001001101111	;
		random_num_table[167]  <= 32'b	00010000111001011010000000111001	;
		random_num_table[168]  <= 32'b	00011100000111110011001011011111	;
		random_num_table[169]  <= 32'b	00000010000000000010000111010001	;
		random_num_table[170]  <= 32'b	00001010010101111110000111111011	;
		random_num_table[171]  <= 32'b	00001111110010000101010101110011	;
		random_num_table[172]  <= 32'b	00010001001110011001001010110011	;
		random_num_table[173]  <= 32'b	00001101010010111010111100111101	;
		random_num_table[174]  <= 32'b	00010000001001000010110000101100	;
		random_num_table[175]  <= 32'b	00010100011100110001100010101111	;
		random_num_table[176]  <= 32'b	00010100011100100001010101110010	;
		random_num_table[177]  <= 32'b	00010010110000000110110000000100	;
		random_num_table[178]  <= 32'b	00010111010000111101001000000000	;
		random_num_table[179]  <= 32'b	00001100010010011000100001011001	;
		random_num_table[180]  <= 32'b	00011110101110100001110000000000	;
		random_num_table[181]  <= 32'b	00000000100001000101000111111100	;
		random_num_table[182]  <= 32'b	00001100000010110100001010100101	;
		random_num_table[183]  <= 32'b	00001000111101010111101100010100	;
		random_num_table[184]  <= 32'b	00011010001100011010011101110011	;
		random_num_table[185]  <= 32'b	00011100010101110111001101000100	;
		random_num_table[186]  <= 32'b	00001100111010011011001110000000	;
		random_num_table[187]  <= 32'b	00001010011010010001010000110101	;
		random_num_table[188]  <= 32'b	00001101010110111011110001010100	;
		random_num_table[189]  <= 32'b	00001010010010111111111000001010	;
		random_num_table[190]  <= 32'b	00001010101000100000010001011100	;
		random_num_table[191]  <= 32'b	00010100000100100101000000110100	;
		random_num_table[192]  <= 32'b	00011111010111011011011110011010	;
		random_num_table[193]  <= 32'b	00010110010100011011100001000001	;
		random_num_table[194]  <= 32'b	00001001110010001010011010101101	;
		random_num_table[195]  <= 32'b	00000000001100000001011111011110	;
		random_num_table[196]  <= 32'b	00011111110011000011010110101010	;
		random_num_table[197]  <= 32'b	00001001111101010001011100010000	;
		random_num_table[198]  <= 32'b	00011100111001110010001000001100	;
		random_num_table[199]  <= 32'b	00011000011011111111101010110110	;
		random_num_table[200]  <= 32'b	00011100011001001010111100111011	;
		random_num_table[201]  <= 32'b	00010001100100100111010101001111	;
		random_num_table[202]  <= 32'b	00010001011001000111111011111001	;
		random_num_table[203]  <= 32'b	00011110111000000011001001110001	;
		random_num_table[204]  <= 32'b	00001000111100010010100001011001	;
		random_num_table[205]  <= 32'b	00011111001010000111001000011100	;
		random_num_table[206]  <= 32'b	00000010001000111010111110001110	;
		random_num_table[207]  <= 32'b	00000000010001001100101111001011	;
		random_num_table[208]  <= 32'b	00000111111000111110111101001001	;
		random_num_table[209]  <= 32'b	00010010000000111011111011000010	;
		random_num_table[210]  <= 32'b	00010110011000011010110011100101	;
		random_num_table[211]  <= 32'b	00000001000100100000010010010010	;
		random_num_table[212]  <= 32'b	00001011001010000000101011010100	;
		random_num_table[213]  <= 32'b	00010111111001111011111011001110	;
		random_num_table[214]  <= 32'b	00011111100100110100011110101110	;
		random_num_table[215]  <= 32'b	00010001110001001000010111100011	;
		random_num_table[216]  <= 32'b	00010000010111011001000100011000	;
		random_num_table[217]  <= 32'b	00000011010011110001100000101101	;
		random_num_table[218]  <= 32'b	00001110101001101010011010111011	;
		random_num_table[219]  <= 32'b	00010101010001000101000010111111	;
		random_num_table[220]  <= 32'b	00010101101111110001000100011110	;
		random_num_table[221]  <= 32'b	00011010111010101010111001010110	;
		random_num_table[222]  <= 32'b	00000110111010111010111000010110	;
		random_num_table[223]  <= 32'b	00011000110111010111000110010011	;
		random_num_table[224]  <= 32'b	00010000100110110010111101000101	;
		random_num_table[225]  <= 32'b	00000010000111000011110000000110	;
		random_num_table[226]  <= 32'b	00001111100011011110001000001000	;
		random_num_table[227]  <= 32'b	00001101010011011001110000101010	;
		random_num_table[228]  <= 32'b	00001000010101011110000000011011	;
		random_num_table[229]  <= 32'b	00001011110101101101010110001011	;
		random_num_table[230]  <= 32'b	00011010011110100111101000001001	;
		random_num_table[231]  <= 32'b	00000000010010111001010110110010	;
		random_num_table[232]  <= 32'b	00001001010001100110000001000101	;
		random_num_table[233]  <= 32'b	00000100111110010100111010100100	;
		random_num_table[234]  <= 32'b	00010001010011011011001010011101	;
		random_num_table[235]  <= 32'b	00001110010011010111100010101011	;
		random_num_table[236]  <= 32'b	00011000000100000110111001011010	;
		random_num_table[237]  <= 32'b	00011111000011111101101100000001	;
		random_num_table[238]  <= 32'b	00011100010010001100001001111010	;
		random_num_table[239]  <= 32'b	00000110111001101001110010100100	;
		random_num_table[240]  <= 32'b	00000110101010001100101100100001	;
		random_num_table[241]  <= 32'b	00000001010000000011001000001110	;
		random_num_table[242]  <= 32'b	00010101001100101110001110111010	;
		random_num_table[243]  <= 32'b	00001001110010000111010001101100	;
		random_num_table[244]  <= 32'b	00001011000111111101100010100110	;
		random_num_table[245]  <= 32'b	00010100110100110010001101111100	;
		random_num_table[246]  <= 32'b	00000110010111101001101011010110	;
		random_num_table[247]  <= 32'b	00000110110110001100100010111010	;
		random_num_table[248]  <= 32'b	00000000010011011001110100110111	;
		random_num_table[249]  <= 32'b	00010110001000110111101011001100	;
		random_num_table[250]  <= 32'b	00001011110110111100100100001010	;
		random_num_table[251]  <= 32'b	00011000111100010110001001011000	;
		random_num_table[252]  <= 32'b	00010000010010000001110001011111	;
		random_num_table[253]  <= 32'b	00000001010100111111110000101011	;
		random_num_table[254]  <= 32'b	00001011001001100000000011110001	;
		random_num_table[255]  <= 32'b	00010001111110101111111110110110	;
	end
endmodule
