`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:54:25 01/19/2015 
// Design Name: 
// Module Name:    rand_table_4 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module rand_table_4(axi_aclk , axi_aresetn , index_num , rand_out , en);
	input			axi_aclk , axi_aresetn , en;
	input		[7:0]	index_num;
	output		[31:0]	rand_out;

	reg 		[31:0]	random_num_table  [255:0];

	assign rand_out = en?random_num_table[index_num]:32'd0;
	
	always@(posedge axi_aclk)
	begin
		random_num_table[0]  <= 32'b	00011010010000001010111000011010	;
		random_num_table[1]  <= 32'b	00011101101010100001001000111001	;
		random_num_table[2]  <= 32'b	00011010100110000111001110111001	;
		random_num_table[3]  <= 32'b	00001101010011100011011111101111	;
		random_num_table[4]  <= 32'b	00011011011100110110101110110001	;
		random_num_table[5]  <= 32'b	00001011101011011100110011010100	;
		random_num_table[6]  <= 32'b	00010101101100110001111110011011	;
		random_num_table[7]  <= 32'b	00011100011010011001010110101101	;
		random_num_table[8]  <= 32'b	00010010001001001111100001110110	;
		random_num_table[9]  <= 32'b	00010001110001010100100101111011	;
		random_num_table[10]  <= 32'b	00001001000110101101100001001010	;
		random_num_table[11]  <= 32'b	00010011010011111001011110000100	;
		random_num_table[12]  <= 32'b	00001000000100101100101100000100	;
		random_num_table[13]  <= 32'b	00001001010111000100000111010001	;
		random_num_table[14]  <= 32'b	00001100001000110010101100100001	;
		random_num_table[15]  <= 32'b	00001000001011000000011001101110	;
		random_num_table[16]  <= 32'b	00010001110101101000011110110011	;
		random_num_table[17]  <= 32'b	00001001011101011101001010100111	;
		random_num_table[18]  <= 32'b	00001111111100110001001000011110	;
		random_num_table[19]  <= 32'b	00000010000110100100010110110111	;
		random_num_table[20]  <= 32'b	00000100101000100101111010111010	;
		random_num_table[21]  <= 32'b	00000001100110101001010010001101	;
		random_num_table[22]  <= 32'b	00000001100010101110010000010001	;
		random_num_table[23]  <= 32'b	00000111001001001110100100111110	;
		random_num_table[24]  <= 32'b	00011010110101000101001000100111	;
		random_num_table[25]  <= 32'b	00010110000111101101001110001100	;
		random_num_table[26]  <= 32'b	00010110011111010100010110111010	;
		random_num_table[27]  <= 32'b	00011010011100000111101111100110	;
		random_num_table[28]  <= 32'b	00000010111100100101111100101001	;
		random_num_table[29]  <= 32'b	00010001100011100010010100011110	;
		random_num_table[30]  <= 32'b	00001001101011100010101001100101	;
		random_num_table[31]  <= 32'b	00000111010101000110011110001000	;
		random_num_table[32]  <= 32'b	00000010011110011001101001010100	;
		random_num_table[33]  <= 32'b	00000100010101110011101001110000	;
		random_num_table[34]  <= 32'b	00011010001110000000010101000010	;
		random_num_table[35]  <= 32'b	00011101000011101000110000011111	;
		random_num_table[36]  <= 32'b	00010101000000000001100010100110	;
		random_num_table[37]  <= 32'b	00001000001100101101000110110011	;
		random_num_table[38]  <= 32'b	00001001101000100100111000000001	;
		random_num_table[39]  <= 32'b	00000111011000100001111001100000	;
		random_num_table[40]  <= 32'b	00000010110010101001000010000000	;
		random_num_table[41]  <= 32'b	00000011100000001110111110100111	;
		random_num_table[42]  <= 32'b	00011101010100001001111101000100	;
		random_num_table[43]  <= 32'b	00001111000001000000111010110110	;
		random_num_table[44]  <= 32'b	00011011000111101110011011001111	;
		random_num_table[45]  <= 32'b	00000110111001011111011010110001	;
		random_num_table[46]  <= 32'b	00011100000010100010111110011101	;
		random_num_table[47]  <= 32'b	00010100111101111001110000111110	;
		random_num_table[48]  <= 32'b	00010101101010000111001101001010	;
		random_num_table[49]  <= 32'b	00010011010001111100100001000011	;
		random_num_table[50]  <= 32'b	00010110110110100010110011011111	;
		random_num_table[51]  <= 32'b	00011001000111001110111001010101	;
		random_num_table[52]  <= 32'b	00000000011011101011011010011110	;
		random_num_table[53]  <= 32'b	00010000100101001010100110101000	;
		random_num_table[54]  <= 32'b	00001100111100111100000101010110	;
		random_num_table[55]  <= 32'b	00000001001011000111111100110010	;
		random_num_table[56]  <= 32'b	00001010010011110101110011011110	;
		random_num_table[57]  <= 32'b	00000111011001011001100110000111	;
		random_num_table[58]  <= 32'b	00010100010000001000100001001100	;
		random_num_table[59]  <= 32'b	00000010001011000010101100101011	;
		random_num_table[60]  <= 32'b	00011001101010101001001101011110	;
		random_num_table[61]  <= 32'b	00011000011001111011100101111010	;
		random_num_table[62]  <= 32'b	00001101001001110100101001010010	;
		random_num_table[63]  <= 32'b	00001111111011000100101110110010	;
		random_num_table[64]  <= 32'b	00000011111111011111001010110111	;
		random_num_table[65]  <= 32'b	00001110111100100011110001010111	;
		random_num_table[66]  <= 32'b	00000110000110010010111100101110	;
		random_num_table[67]  <= 32'b	00011010110110010100010011011101	;
		random_num_table[68]  <= 32'b	00000100011011010111010110010110	;
		random_num_table[69]  <= 32'b	00000011010001010010100011101111	;
		random_num_table[70]  <= 32'b	00010111010011001000100011000001	;
		random_num_table[71]  <= 32'b	00001111010001000100011001010111	;
		random_num_table[72]  <= 32'b	00010101100010101101101110001101	;
		random_num_table[73]  <= 32'b	00010001001010001111011010100101	;
		random_num_table[74]  <= 32'b	00000001011010001110100011001010	;
		random_num_table[75]  <= 32'b	00011010100000010010010101101100	;
		random_num_table[76]  <= 32'b	00011100010001111101110010111011	;
		random_num_table[77]  <= 32'b	00001010001000110011101111010000	;
		random_num_table[78]  <= 32'b	00011110101100110110011101101001	;
		random_num_table[79]  <= 32'b	00011110011001011010011100001100	;
		random_num_table[80]  <= 32'b	00001000110010111011111101010000	;
		random_num_table[81]  <= 32'b	00001100101011101010000000000001	;
		random_num_table[82]  <= 32'b	00010110001110000011001000011010	;
		random_num_table[83]  <= 32'b	00010011101011000000010000111110	;
		random_num_table[84]  <= 32'b	00000010100000011000011001011100	;
		random_num_table[85]  <= 32'b	00011001000111110110111001011001	;
		random_num_table[86]  <= 32'b	00011000111110111001111001000110	;
		random_num_table[87]  <= 32'b	00000100111101110101010100010101	;
		random_num_table[88]  <= 32'b	00000010100100101000000000001010	;
		random_num_table[89]  <= 32'b	00010110101110001000110000001110	;
		random_num_table[90]  <= 32'b	00000100110110001111011101100100	;
		random_num_table[91]  <= 32'b	00010111101110101010011001111010	;
		random_num_table[92]  <= 32'b	00010001101010001100101010101101	;
		random_num_table[93]  <= 32'b	00001111111101101011111001101001	;
		random_num_table[94]  <= 32'b	00011110010000000001010010010101	;
		random_num_table[95]  <= 32'b	00000011101001111010110110010111	;
		random_num_table[96]  <= 32'b	00000100001110111011100100010001	;
		random_num_table[97]  <= 32'b	00010111100011101100100011110100	;
		random_num_table[98]  <= 32'b	00000100111100011100111100101011	;
		random_num_table[99]  <= 32'b	00001110111101001111100001110001	;
		random_num_table[100]  <= 32'b	00010111000001001111100001111100	;
		random_num_table[101]  <= 32'b	00001000100100000110111010110110	;
		random_num_table[102]  <= 32'b	00001001101000001111111011100110	;
		random_num_table[103]  <= 32'b	00001011110010000010010110111010	;
		random_num_table[104]  <= 32'b	00010110001100100101010101101110	;
		random_num_table[105]  <= 32'b	00001100001111111100010111010001	;
		random_num_table[106]  <= 32'b	00011000100110001010000010111101	;
		random_num_table[107]  <= 32'b	00000110000010000100100001101110	;
		random_num_table[108]  <= 32'b	00010111010001110000011000100110	;
		random_num_table[109]  <= 32'b	00010001101010111110011111000000	;
		random_num_table[110]  <= 32'b	00010101110001001110110011110100	;
		random_num_table[111]  <= 32'b	00001010000001101110111100011010	;
		random_num_table[112]  <= 32'b	00001110001111100110000110000010	;
		random_num_table[113]  <= 32'b	00000010001111100011100101101000	;
		random_num_table[114]  <= 32'b	00000001101000100000100000110111	;
		random_num_table[115]  <= 32'b	00011111100000011001010011101010	;
		random_num_table[116]  <= 32'b	00001101000000100010000100100101	;
		random_num_table[117]  <= 32'b	00001010011011000101111111001101	;
		random_num_table[118]  <= 32'b	00000000100110010000001110100100	;
		random_num_table[119]  <= 32'b	00010011100101101001001111111101	;
		random_num_table[120]  <= 32'b	00011011101001110010101101000111	;
		random_num_table[121]  <= 32'b	00011111110000110011110110100101	;
		random_num_table[122]  <= 32'b	00010110101001001111101011111011	;
		random_num_table[123]  <= 32'b	00011100000011101011010010001101	;
		random_num_table[124]  <= 32'b	00011011100011000100001101111111	;
		random_num_table[125]  <= 32'b	00011110101010000010110111000011	;
		random_num_table[126]  <= 32'b	00001011001100110100011110110001	;
		random_num_table[127]  <= 32'b	00010010110011000101010110101000	;
		random_num_table[128]  <= 32'b	00000011011010000101100111101110	;
		random_num_table[129]  <= 32'b	00011001101111101001100000000010	;
		random_num_table[130]  <= 32'b	00001001011001001001101111010101	;
		random_num_table[131]  <= 32'b	00001100101011011001000101110000	;
		random_num_table[132]  <= 32'b	00011110001101010100101011011001	;
		random_num_table[133]  <= 32'b	00000001111111000001111010100100	;
		random_num_table[134]  <= 32'b	00011110011111100000100010001111	;
		random_num_table[135]  <= 32'b	00010001010111101100100111011101	;
		random_num_table[136]  <= 32'b	00001011010001000110111100001000	;
		random_num_table[137]  <= 32'b	00001110011001001011101100111011	;
		random_num_table[138]  <= 32'b	00001011011001110111111000111011	;
		random_num_table[139]  <= 32'b	00001001100010001111001001000110	;
		random_num_table[140]  <= 32'b	00011100101001100010001111110101	;
		random_num_table[141]  <= 32'b	00010111000011101110101110010011	;
		random_num_table[142]  <= 32'b	00010000000100010100110010000010	;
		random_num_table[143]  <= 32'b	00000101011101011100001111011111	;
		random_num_table[144]  <= 32'b	00001111011100011011110011000001	;
		random_num_table[145]  <= 32'b	00001101011100001010100001111001	;
		random_num_table[146]  <= 32'b	00001010001110100101111111010010	;
		random_num_table[147]  <= 32'b	00000000001011001110000010111001	;
		random_num_table[148]  <= 32'b	00001111101100111000111000001101	;
		random_num_table[149]  <= 32'b	00001010000000011111000100111101	;
		random_num_table[150]  <= 32'b	00001111010111100111011001100101	;
		random_num_table[151]  <= 32'b	00011101010001001111101100111100	;
		random_num_table[152]  <= 32'b	00011110110111001110110110101111	;
		random_num_table[153]  <= 32'b	00000010101010000101111111000101	;
		random_num_table[154]  <= 32'b	00000100100001111111001011111001	;
		random_num_table[155]  <= 32'b	00000010010000110000110000001011	;
		random_num_table[156]  <= 32'b	00000111001110110010101001111111	;
		random_num_table[157]  <= 32'b	00000001001000010010110001101100	;
		random_num_table[158]  <= 32'b	00001100010001010110010100011100	;
		random_num_table[159]  <= 32'b	00011111000011001000100010101001	;
		random_num_table[160]  <= 32'b	00001011110111110110100011000110	;
		random_num_table[161]  <= 32'b	00000111110011110101111001111011	;
		random_num_table[162]  <= 32'b	00000011011001110101001010101111	;
		random_num_table[163]  <= 32'b	00010101001000000000110100111010	;
		random_num_table[164]  <= 32'b	00011010010011011110100001111001	;
		random_num_table[165]  <= 32'b	00011000000101000010110110100010	;
		random_num_table[166]  <= 32'b	00011000001010111011001001011110	;
		random_num_table[167]  <= 32'b	00010000101100000001000101110001	;
		random_num_table[168]  <= 32'b	00001110110011110010000010001011	;
		random_num_table[169]  <= 32'b	00001001001001110100011110011011	;
		random_num_table[170]  <= 32'b	00000011110101000011100110000001	;
		random_num_table[171]  <= 32'b	00001100001011110101111110110101	;
		random_num_table[172]  <= 32'b	00011110011111000111010000000111	;
		random_num_table[173]  <= 32'b	00001111001100110110111111110111	;
		random_num_table[174]  <= 32'b	00011010100111001101100110010100	;
		random_num_table[175]  <= 32'b	00011011110111100110111000001101	;
		random_num_table[176]  <= 32'b	00000110000000000101101111110011	;
		random_num_table[177]  <= 32'b	00011101100001101110011000101001	;
		random_num_table[178]  <= 32'b	00010110100011101011000101100010	;
		random_num_table[179]  <= 32'b	00000100110110100000110111011011	;
		random_num_table[180]  <= 32'b	00000100001111101011101001001000	;
		random_num_table[181]  <= 32'b	00000011110011111100001101001111	;
		random_num_table[182]  <= 32'b	00000001100100111001010100011001	;
		random_num_table[183]  <= 32'b	00001010010000000010011011010100	;
		random_num_table[184]  <= 32'b	00000101111111001111100100110110	;
		random_num_table[185]  <= 32'b	00010111010011101001101100101100	;
		random_num_table[186]  <= 32'b	00011101001010010011001110111101	;
		random_num_table[187]  <= 32'b	00010101010011100101100101000101	;
		random_num_table[188]  <= 32'b	00001010101001100011010100111100	;
		random_num_table[189]  <= 32'b	00011111010100111001010011000101	;
		random_num_table[190]  <= 32'b	00011101111001110001010000010111	;
		random_num_table[191]  <= 32'b	00001000000111100001000000010010	;
		random_num_table[192]  <= 32'b	00011110111000010010010000101100	;
		random_num_table[193]  <= 32'b	00011110100111111101001001000000	;
		random_num_table[194]  <= 32'b	00010110001000100011011001010011	;
		random_num_table[195]  <= 32'b	00001001110111111111010110101110	;
		random_num_table[196]  <= 32'b	00011100010011000000100100110100	;
		random_num_table[197]  <= 32'b	00010101001101101000110001111110	;
		random_num_table[198]  <= 32'b	00001110000000110100011010100111	;
		random_num_table[199]  <= 32'b	00010001110000000011001001000111	;
		random_num_table[200]  <= 32'b	00000100110101001001101010111100	;
		random_num_table[201]  <= 32'b	00000100011100001101110101110010	;
		random_num_table[202]  <= 32'b	00001001110111110110000010010001	;
		random_num_table[203]  <= 32'b	00011100110111000001110000101111	;
		random_num_table[204]  <= 32'b	00001110110101110110111100111100	;
		random_num_table[205]  <= 32'b	00000101100100011001100100111000	;
		random_num_table[206]  <= 32'b	00011010011000111010010101001000	;
		random_num_table[207]  <= 32'b	00001111000010011101110010001010	;
		random_num_table[208]  <= 32'b	00010011010001101010110110111010	;
		random_num_table[209]  <= 32'b	00000110000111011100010110000011	;
		random_num_table[210]  <= 32'b	00001111011101010000010010111100	;
		random_num_table[211]  <= 32'b	00000010111101001101010101011111	;
		random_num_table[212]  <= 32'b	00011101111110010000111100111001	;
		random_num_table[213]  <= 32'b	00011100111001001110001100101000	;
		random_num_table[214]  <= 32'b	00001011101110010110011101101111	;
		random_num_table[215]  <= 32'b	00010000010011000111001110100011	;
		random_num_table[216]  <= 32'b	00011001111010100000001100100010	;
		random_num_table[217]  <= 32'b	00001101100011111100010100000000	;
		random_num_table[218]  <= 32'b	00010101110100111101000101110110	;
		random_num_table[219]  <= 32'b	00010000000110101000111100001110	;
		random_num_table[220]  <= 32'b	00011100111000001111010111111000	;
		random_num_table[221]  <= 32'b	00001011111100110110110101111110	;
		random_num_table[222]  <= 32'b	00000010001110010110010100001010	;
		random_num_table[223]  <= 32'b	00011110100011101000110001010000	;
		random_num_table[224]  <= 32'b	00010101101111100110110010100101	;
		random_num_table[225]  <= 32'b	00010011111000111000100111101010	;
		random_num_table[226]  <= 32'b	00011111111010001110011001010100	;
		random_num_table[227]  <= 32'b	00000011100100101100001101101111	;
		random_num_table[228]  <= 32'b	00011000111000010001111100110011	;
		random_num_table[229]  <= 32'b	00011111111100010100101000011110	;
		random_num_table[230]  <= 32'b	00010001011011110101010010011010	;
		random_num_table[231]  <= 32'b	00011101100000111110100001011110	;
		random_num_table[232]  <= 32'b	00010000110000101000010111110111	;
		random_num_table[233]  <= 32'b	00000001010101001000010111100110	;
		random_num_table[234]  <= 32'b	00011000001100010001111110110100	;
		random_num_table[235]  <= 32'b	00011001000001100111001001101010	;
		random_num_table[236]  <= 32'b	00001100000110101001011101101010	;
		random_num_table[237]  <= 32'b	00001110110110011100010001110101	;
		random_num_table[238]  <= 32'b	00011101101111001010010110010001	;
		random_num_table[239]  <= 32'b	00011001011100000001110110110010	;
		random_num_table[240]  <= 32'b	00001001110000010011100100111101	;
		random_num_table[241]  <= 32'b	00000000111010110011010101000100	;
		random_num_table[242]  <= 32'b	00000111011100100001100110110000	;
		random_num_table[243]  <= 32'b	00001010100110110100101011001011	;
		random_num_table[244]  <= 32'b	00001000110000101111100011100100	;
		random_num_table[245]  <= 32'b	00010010001110010110010110111001	;
		random_num_table[246]  <= 32'b	00010011101011110110010100101011	;
		random_num_table[247]  <= 32'b	00011110110111111010111011100111	;
		random_num_table[248]  <= 32'b	00010111111000011011010110101111	;
		random_num_table[249]  <= 32'b	00010011000000010111101110011111	;
		random_num_table[250]  <= 32'b	00010111011011101001001000010111	;
		random_num_table[251]  <= 32'b	00011000100110111101001000100000	;
		random_num_table[252]  <= 32'b	00011110001101001100100110110010	;
		random_num_table[253]  <= 32'b	00011110111001110010101101011111	;
		random_num_table[254]  <= 32'b	00011000110101001000000011011100	;
		random_num_table[255]  <= 32'b	00000010001000110000110010000011	;
	end
endmodule
