`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:32:17 01/18/2015 
// Design Name: 
// Module Name:    rand_table 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module rand_table_0(axi_aclk , axi_aresetn , index_num , rand_out , en);
	input			axi_aclk , axi_aresetn , en;
	input		[7:0]	index_num;
	output		[31:0]	rand_out;

	reg 		[31:0]	random_num_table  [255:0];

	assign rand_out = en?random_num_table[index_num]:32'd0;
	
	always@(posedge axi_aclk)
	begin
		random_num_table[0]  <= 32'b	00010110100110000011000111011100	;
		random_num_table[1]  <= 32'b	00000111111011110110000110001001	;
		random_num_table[2]  <= 32'b	00001011001101110101010111100000	;
		random_num_table[3]  <= 32'b	00001101101011001011101100101101	;
		random_num_table[4]  <= 32'b	00000110100010101011100100111110	;
		random_num_table[5]  <= 32'b	00011100110001100100010111111100	;
		random_num_table[6]  <= 32'b	00001101010000101011001110100110	;
		random_num_table[7]  <= 32'b	00000000011100101001010011101110	;
		random_num_table[8]  <= 32'b	00000111010100110010111001110011	;
		random_num_table[9]  <= 32'b	00001000010010001010001010101011	;
		random_num_table[10]  <= 32'b	00010111101001111100110111100101	;
		random_num_table[11]  <= 32'b	00000110000100101011000101010000	;
		random_num_table[12]  <= 32'b	00011011111111010110000000100000	;
		random_num_table[13]  <= 32'b	00010110010001101110111110100010	;
		random_num_table[14]  <= 32'b	00000110111110111000100000101000	;
		random_num_table[15]  <= 32'b	00011010010001000111001011110010	;
		random_num_table[16]  <= 32'b	00011011111110010101111011110001	;
		random_num_table[17]  <= 32'b	00011010011010110110101111101110	;
		random_num_table[18]  <= 32'b	00011010000100101000111100000111	;
		random_num_table[19]  <= 32'b	00000001011111111011111011101110	;
		random_num_table[20]  <= 32'b	00001010001000100000010000110111	;
		random_num_table[21]  <= 32'b	00011011100110111101110011101101	;
		random_num_table[22]  <= 32'b	00011110001100101110101101011101	;
		random_num_table[23]  <= 32'b	00000001011000011111111110101111	;
		random_num_table[24]  <= 32'b	00000001111010011111110111111010	;
		random_num_table[25]  <= 32'b	00011010101101011100100100110100	;
		random_num_table[26]  <= 32'b	00000000110010110011011010110101	;
		random_num_table[27]  <= 32'b	00001010111111101101100100110110	;
		random_num_table[28]  <= 32'b	00010101000111110010101110100101	;
		random_num_table[29]  <= 32'b	00001011111100101010011001110101	;
		random_num_table[30]  <= 32'b	00000111001100101101110000111110	;
		random_num_table[31]  <= 32'b	00000000000111101110011001011010	;
		random_num_table[32]  <= 32'b	00010011100001101011011101110011	;
		random_num_table[33]  <= 32'b	00000011011000111100101110110000	;
		random_num_table[34]  <= 32'b	00001011001101011100101001010111	;
		random_num_table[35]  <= 32'b	00001100000001000010000000111010	;
		random_num_table[36]  <= 32'b	00001001000011000101100101111111	;
		random_num_table[37]  <= 32'b	00001001101101100100011000011010	;
		random_num_table[38]  <= 32'b	00000101011001011001111010010111	;
		random_num_table[39]  <= 32'b	00001100100111010011010001111100	;
		random_num_table[40]  <= 32'b	00011001100100111100000110011110	;
		random_num_table[41]  <= 32'b	00010011010011111111100001001000	;
		random_num_table[42]  <= 32'b	00001100100001111011101100110011	;
		random_num_table[43]  <= 32'b	00011111100111110011011110010010	;
		random_num_table[44]  <= 32'b	00011100100001000100011111001110	;
		random_num_table[45]  <= 32'b	00000010101100100111000110110010	;
		random_num_table[46]  <= 32'b	00011010111100110001011100010001	;
		random_num_table[47]  <= 32'b	00000110101011001100110001101100	;
		random_num_table[48]  <= 32'b	00001101111011100101001000111011	;
		random_num_table[49]  <= 32'b	00001111010101110010000100100100	;
		random_num_table[50]  <= 32'b	00000100010101000101100000001001	;
		random_num_table[51]  <= 32'b	00010101000000001010010010100101	;
		random_num_table[52]  <= 32'b	00010010000001011010111001101001	;
		random_num_table[53]  <= 32'b	00010101010111001100101001000111	;
		random_num_table[54]  <= 32'b	00001010000100111001100100011111	;
		random_num_table[55]  <= 32'b	00000111101000100111111110100111	;
		random_num_table[56]  <= 32'b	00000000101101111011101101110001	;
		random_num_table[57]  <= 32'b	00011111000011011010000010000001	;
		random_num_table[58]  <= 32'b	00000110001110010101101101111010	;
		random_num_table[59]  <= 32'b	00010001001011011100110010101100	;
		random_num_table[60]  <= 32'b	00000010111100011000110011101001	;
		random_num_table[61]  <= 32'b	00011011101010110000001011000101	;
		random_num_table[62]  <= 32'b	00010001011101111101001101101100	;
		random_num_table[63]  <= 32'b	00000000110111110100111100001100	;
		random_num_table[64]  <= 32'b	00010110111000100001011100110010	;
		random_num_table[65]  <= 32'b	00011010101001101111010101101010	;
		random_num_table[66]  <= 32'b	00010000001111001101001001101000	;
		random_num_table[67]  <= 32'b	00000110100110100010001000111011	;
		random_num_table[68]  <= 32'b	00011111000010100000100110100101	;
		random_num_table[69]  <= 32'b	00000110000000011111000101101010	;
		random_num_table[70]  <= 32'b	00010000000100111011010110011000	;
		random_num_table[71]  <= 32'b	00000011011001110001010001011000	;
		random_num_table[72]  <= 32'b	00011011011110111010000001100111	;
		random_num_table[73]  <= 32'b	00010101001000001111110010011111	;
		random_num_table[74]  <= 32'b	00011101101111010101000110001110	;
		random_num_table[75]  <= 32'b	00010001110100101111000000100111	;
		random_num_table[76]  <= 32'b	00011110010011110010000101111111	;
		random_num_table[77]  <= 32'b	00001011010000111100100100001110	;
		random_num_table[78]  <= 32'b	00011011001010101010010000010101	;
		random_num_table[79]  <= 32'b	00001011110000001111011001001010	;
		random_num_table[80]  <= 32'b	00010101110100110111001011110001	;
		random_num_table[81]  <= 32'b	00010000000101001011010010111011	;
		random_num_table[82]  <= 32'b	00010100011111000110110100001111	;
		random_num_table[83]  <= 32'b	00011011010000001001001011011000	;
		random_num_table[84]  <= 32'b	00010100011110100011111101010010	;
		random_num_table[85]  <= 32'b	00011000101001001011011010011011	;
		random_num_table[86]  <= 32'b	00000000111101010101011000100001	;
		random_num_table[87]  <= 32'b	00010110100001010100100100011000	;
		random_num_table[88]  <= 32'b	00011000110001000011001010111111	;
		random_num_table[89]  <= 32'b	00000010010110111001000011100011	;
		random_num_table[90]  <= 32'b	00010101100011101111011001111011	;
		random_num_table[91]  <= 32'b	00010111000011001111111000001000	;
		random_num_table[92]  <= 32'b	00000110110101001011011101011100	;
		random_num_table[93]  <= 32'b	00011001010001010111001100100111	;
		random_num_table[94]  <= 32'b	00001100001101101001110100110010	;
		random_num_table[95]  <= 32'b	00011010100011001111110010001111	;
		random_num_table[96]  <= 32'b	00001100010111000010101011100011	;
		random_num_table[97]  <= 32'b	00011011010100010111001001110101	;
		random_num_table[98]  <= 32'b	00011110101011010001010001010110	;
		random_num_table[99]  <= 32'b	00001011001110000110011000010100	;
		random_num_table[100]  <= 32'b	00001101111011100101101011001110	;
		random_num_table[101]  <= 32'b	00000001000010001001000011101010	;
		random_num_table[102]  <= 32'b	00000011110000000010000001111110	;
		random_num_table[103]  <= 32'b	00001011110010111111001101101110	;
		random_num_table[104]  <= 32'b	00010111011011000110101000000011	;
		random_num_table[105]  <= 32'b	00000111110000110111110011100101	;
		random_num_table[106]  <= 32'b	00010100110000011100001101000011	;
		random_num_table[107]  <= 32'b	00000111111111001101010111101111	;
		random_num_table[108]  <= 32'b	00011101010110011100011000000010	;
		random_num_table[109]  <= 32'b	00011011001010001100010101100110	;
		random_num_table[110]  <= 32'b	00011100100010000110100100000111	;
		random_num_table[111]  <= 32'b	00001100010110001011001000000110	;
		random_num_table[112]  <= 32'b	00011100001111000010000010110011	;
		random_num_table[113]  <= 32'b	00001111110111011000001010100100	;
		random_num_table[114]  <= 32'b	00011111110000010010110111010111	;
		random_num_table[115]  <= 32'b	00001000111000010010000001011011	;
		random_num_table[116]  <= 32'b	00000011001001001110001001010001	;
		random_num_table[117]  <= 32'b	00011110101110011101011111000000	;
		random_num_table[118]  <= 32'b	00001111010111110000010001100001	;
		random_num_table[119]  <= 32'b	00011001110100101110011010001011	;
		random_num_table[120]  <= 32'b	00000111000010100101011011110001	;
		random_num_table[121]  <= 32'b	00011000110111001110110101010001	;
		random_num_table[122]  <= 32'b	00000001101110010101101110010101	;
		random_num_table[123]  <= 32'b	00000111110011001111100001100001	;
		random_num_table[124]  <= 32'b	00010101110111101101001111000101	;
		random_num_table[125]  <= 32'b	00010110100001111000001011001110	;
		random_num_table[126]  <= 32'b	00010001101100101000010110110100	;
		random_num_table[127]  <= 32'b	00001100001011000011010110011100	;
		random_num_table[128]  <= 32'b	00000110111000101100001111111001	;
		random_num_table[129]  <= 32'b	00001111000110100111010010100011	;
		random_num_table[130]  <= 32'b	00001011001000011010101101010011	;
		random_num_table[131]  <= 32'b	00001111001010011110111000110100	;
		random_num_table[132]  <= 32'b	00000001010101001100110110010000	;
		random_num_table[133]  <= 32'b	00011101001001000101110111011100	;
		random_num_table[134]  <= 32'b	00000111110011101111001001010010	;
		random_num_table[135]  <= 32'b	00011111000110101000011001111000	;
		random_num_table[136]  <= 32'b	00010010100111110100011011111110	;
		random_num_table[137]  <= 32'b	00000010011101010011111101110110	;
		random_num_table[138]  <= 32'b	00000001010100110001000001011110	;
		random_num_table[139]  <= 32'b	00011111001100110010000010100010	;
		random_num_table[140]  <= 32'b	00001111110001100100010001101011	;
		random_num_table[141]  <= 32'b	00001101111011100110000110100110	;
		random_num_table[142]  <= 32'b	00001111011101110101101101101110	;
		random_num_table[143]  <= 32'b	00010000010100001111101111011111	;
		random_num_table[144]  <= 32'b	00011110110100011001100010111000	;
		random_num_table[145]  <= 32'b	00010100001001000011000101001000	;
		random_num_table[146]  <= 32'b	00000111000000110000000000010001	;
		random_num_table[147]  <= 32'b	00010010001100010001010111000101	;
		random_num_table[148]  <= 32'b	00000001101000010100100000011000	;
		random_num_table[149]  <= 32'b	00010001011001001110111001011111	;
		random_num_table[150]  <= 32'b	00001001010001101000101000100111	;
		random_num_table[151]  <= 32'b	00000001110110001100111010111011	;
		random_num_table[152]  <= 32'b	00010001001110011000100101110110	;
		random_num_table[153]  <= 32'b	00001010100110000010101110110010	;
		random_num_table[154]  <= 32'b	00011100111110011011010110000011	;
		random_num_table[155]  <= 32'b	00001101101100010111001101101101	;
		random_num_table[156]  <= 32'b	00001011110000111111110000001101	;
		random_num_table[157]  <= 32'b	00010001110110101110000100101100	;
		random_num_table[158]  <= 32'b	00011010101011111100001100100001	;
		random_num_table[159]  <= 32'b	00000010010011111000001000111001	;
		random_num_table[160]  <= 32'b	00011111011010010000111010101111	;
		random_num_table[161]  <= 32'b	00001100010111111101101110110001	;
		random_num_table[162]  <= 32'b	00010011000011011010110111001110	;
		random_num_table[163]  <= 32'b	00011010010101110001011101010101	;
		random_num_table[164]  <= 32'b	00011011010110011101011001011010	;
		random_num_table[165]  <= 32'b	00010010110100011000001110001111	;
		random_num_table[166]  <= 32'b	00001110011110101000111100000111	;
		random_num_table[167]  <= 32'b	00001111000100001011100100001110	;
		random_num_table[168]  <= 32'b	00011010111101111010010010111100	;
		random_num_table[169]  <= 32'b	00001011001100100001100011111110	;
		random_num_table[170]  <= 32'b	00000101110001100000111111001101	;
		random_num_table[171]  <= 32'b	00010111111101000100100100000110	;
		random_num_table[172]  <= 32'b	00000111001101101111111101100001	;
		random_num_table[173]  <= 32'b	00000000010000100011100110101111	;
		random_num_table[174]  <= 32'b	00011111101001000101011010100110	;
		random_num_table[175]  <= 32'b	00011011101010100011000100111101	;
		random_num_table[176]  <= 32'b	00010000001111111111100101000110	;
		random_num_table[177]  <= 32'b	00011101101110000110001110001101	;
		random_num_table[178]  <= 32'b	00010000111000100100001101101000	;
		random_num_table[179]  <= 32'b	00011011100111111001100011101100	;
		random_num_table[180]  <= 32'b	00001100111110101010011000011100	;
		random_num_table[181]  <= 32'b	00010001000000010000111111011100	;
		random_num_table[182]  <= 32'b	00001110101000110011100111011101	;
		random_num_table[183]  <= 32'b	00001101001110000100110000100110	;
		random_num_table[184]  <= 32'b	00000110110110010000111011100101	;
		random_num_table[185]  <= 32'b	00010010101110101100110100010111	;
		random_num_table[186]  <= 32'b	00000010100111011101110101011001	;
		random_num_table[187]  <= 32'b	00001010110101100011101100001001	;
		random_num_table[188]  <= 32'b	00001010010101101111011101100000	;
		random_num_table[189]  <= 32'b	00011010010011100010100101011101	;
		random_num_table[190]  <= 32'b	00010111001000000000011011100110	;
		random_num_table[191]  <= 32'b	00000001001010011111001000011100	;
		random_num_table[192]  <= 32'b	00000001001011010100100011111101	;
		random_num_table[193]  <= 32'b	00011100101011100010011011100110	;
		random_num_table[194]  <= 32'b	00011000101110011010111110101101	;
		random_num_table[195]  <= 32'b	00001000101000100001011111111001	;
		random_num_table[196]  <= 32'b	00011000110010101001000011010111	;
		random_num_table[197]  <= 32'b	00011100000010001110101111001111	;
		random_num_table[198]  <= 32'b	00011101101101101110010111010011	;
		random_num_table[199]  <= 32'b	00000111100000000000010011001110	;
		random_num_table[200]  <= 32'b	00011000011000011001110000110111	;
		random_num_table[201]  <= 32'b	00010000101001011000100101010001	;
		random_num_table[202]  <= 32'b	00010010110100110011110011011001	;
		random_num_table[203]  <= 32'b	00000010100111001100100101010000	;
		random_num_table[204]  <= 32'b	00000111101111101100001100000110	;
		random_num_table[205]  <= 32'b	00000111100001000001100110100101	;
		random_num_table[206]  <= 32'b	00001101100111011110110111010011	;
		random_num_table[207]  <= 32'b	00000000001000001000100011111000	;
		random_num_table[208]  <= 32'b	00000111010000111100011101101110	;
		random_num_table[209]  <= 32'b	00010010111111010011111110000011	;
		random_num_table[210]  <= 32'b	00010111110000001101001101011011	;
		random_num_table[211]  <= 32'b	00001001011100011110000110111110	;
		random_num_table[212]  <= 32'b	00001101101110010000011011000011	;
		random_num_table[213]  <= 32'b	00011100010010111100010101101001	;
		random_num_table[214]  <= 32'b	00010111010100100101001000000101	;
		random_num_table[215]  <= 32'b	00010101001001011001010000110011	;
		random_num_table[216]  <= 32'b	00000101111000110110001111000000	;
		random_num_table[217]  <= 32'b	00010011100011000011000000011101	;
		random_num_table[218]  <= 32'b	00001001110010111000000000101111	;
		random_num_table[219]  <= 32'b	00010100000111000110101101011100	;
		random_num_table[220]  <= 32'b	00011111010011011000100001110100	;
		random_num_table[221]  <= 32'b	00000110111010101000010110001011	;
		random_num_table[222]  <= 32'b	00010101000010110101010001101101	;
		random_num_table[223]  <= 32'b	00011100010100111001100000011000	;
		random_num_table[224]  <= 32'b	00000101111010011111101011110101	;
		random_num_table[225]  <= 32'b	00001000111111011110111010011001	;
		random_num_table[226]  <= 32'b	00010110110001111111111100000010	;
		random_num_table[227]  <= 32'b	00011011011001111111010110011001	;
		random_num_table[228]  <= 32'b	00000100001001010000110110110001	;
		random_num_table[229]  <= 32'b	00001100001111100100001010001111	;
		random_num_table[230]  <= 32'b	00011110011000111110110011110110	;
		random_num_table[231]  <= 32'b	00010011010010110110100110011000	;
		random_num_table[232]  <= 32'b	00000100001001000010111010111010	;
		random_num_table[233]  <= 32'b	00011100010110011011011110011110	;
		random_num_table[234]  <= 32'b	00011011101001000010010111010000	;
		random_num_table[235]  <= 32'b	00000011001100100011001000001110	;
		random_num_table[236]  <= 32'b	00001001101100101010111100111110	;
		random_num_table[237]  <= 32'b	00000101011110111100000111011000	;
		random_num_table[238]  <= 32'b	00000000110010101110101100011001	;
		random_num_table[239]  <= 32'b	00010101111010011100010010000110	;
		random_num_table[240]  <= 32'b	00001101101011000111011101001110	;
		random_num_table[241]  <= 32'b	00001101000011110101010100011101	;
		random_num_table[242]  <= 32'b	00010111000100110101110100010110	;
		random_num_table[243]  <= 32'b	00000100101101011000010111011010	;
		random_num_table[244]  <= 32'b	00001001110011110111010011101011	;
		random_num_table[245]  <= 32'b	00010110000011000011101111100000	;
		random_num_table[246]  <= 32'b	00010001010110100010100011110010	;
		random_num_table[247]  <= 32'b	00001001000001101001001110110011	;
		random_num_table[248]  <= 32'b	00001100100001010000011001011110	;
		random_num_table[249]  <= 32'b	00010100011100100001000000001011	;
		random_num_table[250]  <= 32'b	00001010010010000111110101111011	;
		random_num_table[251]  <= 32'b	00010101000101101000011101001011	;
		random_num_table[252]  <= 32'b	00001110010101000101110001001000	;
		random_num_table[253]  <= 32'b	00011000010100111111011001010111	;
		random_num_table[254]  <= 32'b	00011011000010111110011110010010	;
		random_num_table[255]  <= 32'b	00011100011010111110101000111100	;
	end

endmodule
