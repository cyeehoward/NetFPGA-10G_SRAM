`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:20:22 02/01/2016 
// Design Name: 
// Module Name:    packet_collector 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module packet_collector(inc , inc_tuser , sum_tdata , sum_tdata_valid , sum_tuser , sum_tuser_valid , memclk , reset , tuser , dout_valid_tuser , axififo_din , axififo_din_valid , axififo_empty , rempty_tuser , axififo_mem_queue_full);
	input																memclk , reset;	
	input  															axififo_empty;
	input  	[((8*24+9)-1):0]			axififo_din;	
	input  	        												axififo_din_valid;
	input 	[(128 - 1):0] 							tuser;
	input 	 														dout_valid_tuser;
	input 	 														rempty_tuser;
	input 			        										axififo_mem_queue_full;
	output reg 														inc;
	output reg 														inc_tuser;
	output reg   	[((8*24+9)-1):0]	sum_tdata;	
	output reg  	[(128 - 1):0] 		sum_tuser;
	output reg   							sum_tdata_valid;	
	output reg  							sum_tuser_valid;
	////////////////////////////////////////////////////////////////
	//save packet 
	reg	[200:0]				tdata_save	[255:0];
   reg 	[127:0]          	tuser_save		[255:0];
	reg	[1:0]					count_clk;
	reg	[1:0]					count_packet;
	reg	[8:0]		packet_num_count;
	////////////////////////////////////////////////////////////////	
	reg	[15:0]				eth_type;
	always@(*)
	begin
		if(axififo_din_valid)
		begin
			eth_type[15:8]	= axififo_din[112:105];
			eth_type[7:0]	= axififo_din[120:113];	
		end
		else
		begin
			eth_type 		= 16'd0;
		end
	end
	////////////////////////////////////////////////////////////////
	
	always@(posedge memclk or negedge reset)
	begin
		if(~reset)
		begin
			tdata_save	[	0	]	<=	201'd0	;
			tdata_save	[	1	]	<=	201'd0	;
			tdata_save	[	2	]	<=	201'd0	;
			tdata_save	[	3	]	<=	201'd0	;
			tdata_save	[	4	]	<=	201'd0	;
			tdata_save	[	5	]	<=	201'd0	;
			tdata_save	[	6	]	<=	201'd0	;
			tdata_save	[	7	]	<=	201'd0	;
			tdata_save	[	8	]	<=	201'd0	;
			tdata_save	[	9	]	<=	201'd0	;
			tdata_save	[	10	]	<=	201'd0	;
			tdata_save	[	11	]	<=	201'd0	;
			tdata_save	[	12	]	<=	201'd0	;
			tdata_save	[	13	]	<=	201'd0	;
			tdata_save	[	14	]	<=	201'd0	;
			tdata_save	[	15	]	<=	201'd0	;
			tdata_save	[	16	]	<=	201'd0	;
			tdata_save	[	17	]	<=	201'd0	;
			tdata_save	[	18	]	<=	201'd0	;
			tdata_save	[	19	]	<=	201'd0	;
			tdata_save	[	20	]	<=	201'd0	;
			tdata_save	[	21	]	<=	201'd0	;
			tdata_save	[	22	]	<=	201'd0	;
			tdata_save	[	23	]	<=	201'd0	;
			tdata_save	[	24	]	<=	201'd0	;
			tdata_save	[	25	]	<=	201'd0	;
			tdata_save	[	26	]	<=	201'd0	;
			tdata_save	[	27	]	<=	201'd0	;
			tdata_save	[	28	]	<=	201'd0	;
			tdata_save	[	29	]	<=	201'd0	;
			tdata_save	[	30	]	<=	201'd0	;
			tdata_save	[	31	]	<=	201'd0	;
			tdata_save	[	32	]	<=	201'd0	;
			tdata_save	[	33	]	<=	201'd0	;
			tdata_save	[	34	]	<=	201'd0	;
			tdata_save	[	35	]	<=	201'd0	;
			tdata_save	[	36	]	<=	201'd0	;
			tdata_save	[	37	]	<=	201'd0	;
			tdata_save	[	38	]	<=	201'd0	;
			tdata_save	[	39	]	<=	201'd0	;
			tdata_save	[	40	]	<=	201'd0	;
			tdata_save	[	41	]	<=	201'd0	;
			tdata_save	[	42	]	<=	201'd0	;
			tdata_save	[	43	]	<=	201'd0	;
			tdata_save	[	44	]	<=	201'd0	;
			tdata_save	[	45	]	<=	201'd0	;
			tdata_save	[	46	]	<=	201'd0	;
			tdata_save	[	47	]	<=	201'd0	;
			tdata_save	[	48	]	<=	201'd0	;
			tdata_save	[	49	]	<=	201'd0	;
			tdata_save	[	50	]	<=	201'd0	;
			tdata_save	[	51	]	<=	201'd0	;
			tdata_save	[	52	]	<=	201'd0	;
			tdata_save	[	53	]	<=	201'd0	;
			tdata_save	[	54	]	<=	201'd0	;
			tdata_save	[	55	]	<=	201'd0	;
			tdata_save	[	56	]	<=	201'd0	;
			tdata_save	[	57	]	<=	201'd0	;
			tdata_save	[	58	]	<=	201'd0	;
			tdata_save	[	59	]	<=	201'd0	;
			tdata_save	[	60	]	<=	201'd0	;
			tdata_save	[	61	]	<=	201'd0	;
			tdata_save	[	62	]	<=	201'd0	;
			tdata_save	[	63	]	<=	201'd0	;
			tdata_save	[	64	]	<=	201'd0	;
			tdata_save	[	65	]	<=	201'd0	;
			tdata_save	[	66	]	<=	201'd0	;
			tdata_save	[	67	]	<=	201'd0	;
			tdata_save	[	68	]	<=	201'd0	;
			tdata_save	[	69	]	<=	201'd0	;
			tdata_save	[	70	]	<=	201'd0	;
			tdata_save	[	71	]	<=	201'd0	;
			tdata_save	[	72	]	<=	201'd0	;
			tdata_save	[	73	]	<=	201'd0	;
			tdata_save	[	74	]	<=	201'd0	;
			tdata_save	[	75	]	<=	201'd0	;
			tdata_save	[	76	]	<=	201'd0	;
			tdata_save	[	77	]	<=	201'd0	;
			tdata_save	[	78	]	<=	201'd0	;
			tdata_save	[	79	]	<=	201'd0	;
			tdata_save	[	80	]	<=	201'd0	;
			tdata_save	[	81	]	<=	201'd0	;
			tdata_save	[	82	]	<=	201'd0	;
			tdata_save	[	83	]	<=	201'd0	;
			tdata_save	[	84	]	<=	201'd0	;
			tdata_save	[	85	]	<=	201'd0	;
			tdata_save	[	86	]	<=	201'd0	;
			tdata_save	[	87	]	<=	201'd0	;
			tdata_save	[	88	]	<=	201'd0	;
			tdata_save	[	89	]	<=	201'd0	;
			tdata_save	[	90	]	<=	201'd0	;
			tdata_save	[	91	]	<=	201'd0	;
			tdata_save	[	92	]	<=	201'd0	;
			tdata_save	[	93	]	<=	201'd0	;
			tdata_save	[	94	]	<=	201'd0	;
			tdata_save	[	95	]	<=	201'd0	;
			tdata_save	[	96	]	<=	201'd0	;
			tdata_save	[	97	]	<=	201'd0	;
			tdata_save	[	98	]	<=	201'd0	;
			tdata_save	[	99	]	<=	201'd0	;
			tdata_save	[	100	]	<=	201'd0	;
			tdata_save	[	101	]	<=	201'd0	;
			tdata_save	[	102	]	<=	201'd0	;
			tdata_save	[	103	]	<=	201'd0	;
			tdata_save	[	104	]	<=	201'd0	;
			tdata_save	[	105	]	<=	201'd0	;
			tdata_save	[	106	]	<=	201'd0	;
			tdata_save	[	107	]	<=	201'd0	;
			tdata_save	[	108	]	<=	201'd0	;
			tdata_save	[	109	]	<=	201'd0	;
			tdata_save	[	110	]	<=	201'd0	;
			tdata_save	[	111	]	<=	201'd0	;
			tdata_save	[	112	]	<=	201'd0	;
			tdata_save	[	113	]	<=	201'd0	;
			tdata_save	[	114	]	<=	201'd0	;
			tdata_save	[	115	]	<=	201'd0	;
			tdata_save	[	116	]	<=	201'd0	;
			tdata_save	[	117	]	<=	201'd0	;
			tdata_save	[	118	]	<=	201'd0	;
			tdata_save	[	119	]	<=	201'd0	;
			tdata_save	[	120	]	<=	201'd0	;
			tdata_save	[	121	]	<=	201'd0	;
			tdata_save	[	122	]	<=	201'd0	;
			tdata_save	[	123	]	<=	201'd0	;
			tdata_save	[	124	]	<=	201'd0	;
			tdata_save	[	125	]	<=	201'd0	;
			tdata_save	[	126	]	<=	201'd0	;
			tdata_save	[	127	]	<=	201'd0	;
			tdata_save	[	128	]	<=	201'd0	;
			tdata_save	[	129	]	<=	201'd0	;
			tdata_save	[	130	]	<=	201'd0	;
			tdata_save	[	131	]	<=	201'd0	;
			tdata_save	[	132	]	<=	201'd0	;
			tdata_save	[	133	]	<=	201'd0	;
			tdata_save	[	134	]	<=	201'd0	;
			tdata_save	[	135	]	<=	201'd0	;
			tdata_save	[	136	]	<=	201'd0	;
			tdata_save	[	137	]	<=	201'd0	;
			tdata_save	[	138	]	<=	201'd0	;
			tdata_save	[	139	]	<=	201'd0	;
			tdata_save	[	140	]	<=	201'd0	;
			tdata_save	[	141	]	<=	201'd0	;
			tdata_save	[	142	]	<=	201'd0	;
			tdata_save	[	143	]	<=	201'd0	;
			tdata_save	[	144	]	<=	201'd0	;
			tdata_save	[	145	]	<=	201'd0	;
			tdata_save	[	146	]	<=	201'd0	;
			tdata_save	[	147	]	<=	201'd0	;
			tdata_save	[	148	]	<=	201'd0	;
			tdata_save	[	149	]	<=	201'd0	;
			tdata_save	[	150	]	<=	201'd0	;
			tdata_save	[	151	]	<=	201'd0	;
			tdata_save	[	152	]	<=	201'd0	;
			tdata_save	[	153	]	<=	201'd0	;
			tdata_save	[	154	]	<=	201'd0	;
			tdata_save	[	155	]	<=	201'd0	;
			tdata_save	[	156	]	<=	201'd0	;
			tdata_save	[	157	]	<=	201'd0	;
			tdata_save	[	158	]	<=	201'd0	;
			tdata_save	[	159	]	<=	201'd0	;
			tdata_save	[	160	]	<=	201'd0	;
			tdata_save	[	161	]	<=	201'd0	;
			tdata_save	[	162	]	<=	201'd0	;
			tdata_save	[	163	]	<=	201'd0	;
			tdata_save	[	164	]	<=	201'd0	;
			tdata_save	[	165	]	<=	201'd0	;
			tdata_save	[	166	]	<=	201'd0	;
			tdata_save	[	167	]	<=	201'd0	;
			tdata_save	[	168	]	<=	201'd0	;
			tdata_save	[	169	]	<=	201'd0	;
			tdata_save	[	170	]	<=	201'd0	;
			tdata_save	[	171	]	<=	201'd0	;
			tdata_save	[	172	]	<=	201'd0	;
			tdata_save	[	173	]	<=	201'd0	;
			tdata_save	[	174	]	<=	201'd0	;
			tdata_save	[	175	]	<=	201'd0	;
			tdata_save	[	176	]	<=	201'd0	;
			tdata_save	[	177	]	<=	201'd0	;
			tdata_save	[	178	]	<=	201'd0	;
			tdata_save	[	179	]	<=	201'd0	;
			tdata_save	[	180	]	<=	201'd0	;
			tdata_save	[	181	]	<=	201'd0	;
			tdata_save	[	182	]	<=	201'd0	;
			tdata_save	[	183	]	<=	201'd0	;
			tdata_save	[	184	]	<=	201'd0	;
			tdata_save	[	185	]	<=	201'd0	;
			tdata_save	[	186	]	<=	201'd0	;
			tdata_save	[	187	]	<=	201'd0	;
			tdata_save	[	188	]	<=	201'd0	;
			tdata_save	[	189	]	<=	201'd0	;
			tdata_save	[	190	]	<=	201'd0	;
			tdata_save	[	191	]	<=	201'd0	;
			tdata_save	[	192	]	<=	201'd0	;
			tdata_save	[	193	]	<=	201'd0	;
			tdata_save	[	194	]	<=	201'd0	;
			tdata_save	[	195	]	<=	201'd0	;
			tdata_save	[	196	]	<=	201'd0	;
			tdata_save	[	197	]	<=	201'd0	;
			tdata_save	[	198	]	<=	201'd0	;
			tdata_save	[	199	]	<=	201'd0	;
			tdata_save	[	200	]	<=	201'd0	;
			tdata_save	[	201	]	<=	201'd0	;
			tdata_save	[	202	]	<=	201'd0	;
			tdata_save	[	203	]	<=	201'd0	;
			tdata_save	[	204	]	<=	201'd0	;
			tdata_save	[	205	]	<=	201'd0	;
			tdata_save	[	206	]	<=	201'd0	;
			tdata_save	[	207	]	<=	201'd0	;
			tdata_save	[	208	]	<=	201'd0	;
			tdata_save	[	209	]	<=	201'd0	;
			tdata_save	[	210	]	<=	201'd0	;
			tdata_save	[	211	]	<=	201'd0	;
			tdata_save	[	212	]	<=	201'd0	;
			tdata_save	[	213	]	<=	201'd0	;
			tdata_save	[	214	]	<=	201'd0	;
			tdata_save	[	215	]	<=	201'd0	;
			tdata_save	[	216	]	<=	201'd0	;
			tdata_save	[	217	]	<=	201'd0	;
			tdata_save	[	218	]	<=	201'd0	;
			tdata_save	[	219	]	<=	201'd0	;
			tdata_save	[	220	]	<=	201'd0	;
			tdata_save	[	221	]	<=	201'd0	;
			tdata_save	[	222	]	<=	201'd0	;
			tdata_save	[	223	]	<=	201'd0	;
			tdata_save	[	224	]	<=	201'd0	;
			tdata_save	[	225	]	<=	201'd0	;
			tdata_save	[	226	]	<=	201'd0	;
			tdata_save	[	227	]	<=	201'd0	;
			tdata_save	[	228	]	<=	201'd0	;
			tdata_save	[	229	]	<=	201'd0	;
			tdata_save	[	230	]	<=	201'd0	;
			tdata_save	[	231	]	<=	201'd0	;
			tdata_save	[	232	]	<=	201'd0	;
			tdata_save	[	233	]	<=	201'd0	;
			tdata_save	[	234	]	<=	201'd0	;
			tdata_save	[	235	]	<=	201'd0	;
			tdata_save	[	236	]	<=	201'd0	;
			tdata_save	[	237	]	<=	201'd0	;
			tdata_save	[	238	]	<=	201'd0	;
			tdata_save	[	239	]	<=	201'd0	;
			tdata_save	[	240	]	<=	201'd0	;
			tdata_save	[	241	]	<=	201'd0	;
			tdata_save	[	242	]	<=	201'd0	;
			tdata_save	[	243	]	<=	201'd0	;
			tdata_save	[	244	]	<=	201'd0	;
			tdata_save	[	245	]	<=	201'd0	;
			tdata_save	[	246	]	<=	201'd0	;
			tdata_save	[	247	]	<=	201'd0	;
			tdata_save	[	248	]	<=	201'd0	;
			tdata_save	[	249	]	<=	201'd0	;
			tdata_save	[	250	]	<=	201'd0	;
			tdata_save	[	251	]	<=	201'd0	;
			tdata_save	[	252	]	<=	201'd0	;
			tdata_save	[	253	]	<=	201'd0	;
			tdata_save	[	254	]	<=	201'd0	;
			tdata_save	[	255	]	<=	201'd0	;
			tuser_save	[	0	]	<=	128'd0	;
				tuser_save	[	1	]	<=	128'd0	;
				tuser_save	[	2	]	<=	128'd0	;
				tuser_save	[	3	]	<=	128'd0	;
				tuser_save	[	4	]	<=	128'd0	;
				tuser_save	[	5	]	<=	128'd0	;
				tuser_save	[	6	]	<=	128'd0	;
				tuser_save	[	7	]	<=	128'd0	;
				tuser_save	[	8	]	<=	128'd0	;
				tuser_save	[	9	]	<=	128'd0	;
				tuser_save	[	10	]	<=	128'd0	;
				tuser_save	[	11	]	<=	128'd0	;
				tuser_save	[	12	]	<=	128'd0	;
				tuser_save	[	13	]	<=	128'd0	;
				tuser_save	[	14	]	<=	128'd0	;
				tuser_save	[	15	]	<=	128'd0	;
				tuser_save	[	16	]	<=	128'd0	;
				tuser_save	[	17	]	<=	128'd0	;
				tuser_save	[	18	]	<=	128'd0	;
				tuser_save	[	19	]	<=	128'd0	;
				tuser_save	[	20	]	<=	128'd0	;
				tuser_save	[	21	]	<=	128'd0	;
				tuser_save	[	22	]	<=	128'd0	;
				tuser_save	[	23	]	<=	128'd0	;
				tuser_save	[	24	]	<=	128'd0	;
				tuser_save	[	25	]	<=	128'd0	;
				tuser_save	[	26	]	<=	128'd0	;
				tuser_save	[	27	]	<=	128'd0	;
				tuser_save	[	28	]	<=	128'd0	;
				tuser_save	[	29	]	<=	128'd0	;
				tuser_save	[	30	]	<=	128'd0	;
				tuser_save	[	31	]	<=	128'd0	;
				tuser_save	[	32	]	<=	128'd0	;
				tuser_save	[	33	]	<=	128'd0	;
				tuser_save	[	34	]	<=	128'd0	;
				tuser_save	[	35	]	<=	128'd0	;
				tuser_save	[	36	]	<=	128'd0	;
				tuser_save	[	37	]	<=	128'd0	;
				tuser_save	[	38	]	<=	128'd0	;
				tuser_save	[	39	]	<=	128'd0	;
				tuser_save	[	40	]	<=	128'd0	;
				tuser_save	[	41	]	<=	128'd0	;
				tuser_save	[	42	]	<=	128'd0	;
				tuser_save	[	43	]	<=	128'd0	;
				tuser_save	[	44	]	<=	128'd0	;
				tuser_save	[	45	]	<=	128'd0	;
				tuser_save	[	46	]	<=	128'd0	;
				tuser_save	[	47	]	<=	128'd0	;
				tuser_save	[	48	]	<=	128'd0	;
				tuser_save	[	49	]	<=	128'd0	;
				tuser_save	[	50	]	<=	128'd0	;
				tuser_save	[	51	]	<=	128'd0	;
				tuser_save	[	52	]	<=	128'd0	;
				tuser_save	[	53	]	<=	128'd0	;
				tuser_save	[	54	]	<=	128'd0	;
				tuser_save	[	55	]	<=	128'd0	;
				tuser_save	[	56	]	<=	128'd0	;
				tuser_save	[	57	]	<=	128'd0	;
				tuser_save	[	58	]	<=	128'd0	;
				tuser_save	[	59	]	<=	128'd0	;
				tuser_save	[	60	]	<=	128'd0	;
				tuser_save	[	61	]	<=	128'd0	;
				tuser_save	[	62	]	<=	128'd0	;
				tuser_save	[	63	]	<=	128'd0	;
				tuser_save	[	64	]	<=	128'd0	;
				tuser_save	[	65	]	<=	128'd0	;
				tuser_save	[	66	]	<=	128'd0	;
				tuser_save	[	67	]	<=	128'd0	;
				tuser_save	[	68	]	<=	128'd0	;
				tuser_save	[	69	]	<=	128'd0	;
				tuser_save	[	70	]	<=	128'd0	;
				tuser_save	[	71	]	<=	128'd0	;
				tuser_save	[	72	]	<=	128'd0	;
				tuser_save	[	73	]	<=	128'd0	;
				tuser_save	[	74	]	<=	128'd0	;
				tuser_save	[	75	]	<=	128'd0	;
				tuser_save	[	76	]	<=	128'd0	;
				tuser_save	[	77	]	<=	128'd0	;
				tuser_save	[	78	]	<=	128'd0	;
				tuser_save	[	79	]	<=	128'd0	;
				tuser_save	[	80	]	<=	128'd0	;
				tuser_save	[	81	]	<=	128'd0	;
				tuser_save	[	82	]	<=	128'd0	;
				tuser_save	[	83	]	<=	128'd0	;
				tuser_save	[	84	]	<=	128'd0	;
				tuser_save	[	85	]	<=	128'd0	;
				tuser_save	[	86	]	<=	128'd0	;
				tuser_save	[	87	]	<=	128'd0	;
				tuser_save	[	88	]	<=	128'd0	;
				tuser_save	[	89	]	<=	128'd0	;
				tuser_save	[	90	]	<=	128'd0	;
				tuser_save	[	91	]	<=	128'd0	;
				tuser_save	[	92	]	<=	128'd0	;
				tuser_save	[	93	]	<=	128'd0	;
				tuser_save	[	94	]	<=	128'd0	;
				tuser_save	[	95	]	<=	128'd0	;
				tuser_save	[	96	]	<=	128'd0	;
				tuser_save	[	97	]	<=	128'd0	;
				tuser_save	[	98	]	<=	128'd0	;
				tuser_save	[	99	]	<=	128'd0	;
				tuser_save	[	100	]	<=	128'd0	;
				tuser_save	[	101	]	<=	128'd0	;
				tuser_save	[	102	]	<=	128'd0	;
				tuser_save	[	103	]	<=	128'd0	;
				tuser_save	[	104	]	<=	128'd0	;
				tuser_save	[	105	]	<=	128'd0	;
				tuser_save	[	106	]	<=	128'd0	;
				tuser_save	[	107	]	<=	128'd0	;
				tuser_save	[	108	]	<=	128'd0	;
				tuser_save	[	109	]	<=	128'd0	;
				tuser_save	[	110	]	<=	128'd0	;
				tuser_save	[	111	]	<=	128'd0	;
				tuser_save	[	112	]	<=	128'd0	;
				tuser_save	[	113	]	<=	128'd0	;
				tuser_save	[	114	]	<=	128'd0	;
				tuser_save	[	115	]	<=	128'd0	;
				tuser_save	[	116	]	<=	128'd0	;
				tuser_save	[	117	]	<=	128'd0	;
				tuser_save	[	118	]	<=	128'd0	;
				tuser_save	[	119	]	<=	128'd0	;
				tuser_save	[	120	]	<=	128'd0	;
				tuser_save	[	121	]	<=	128'd0	;
				tuser_save	[	122	]	<=	128'd0	;
				tuser_save	[	123	]	<=	128'd0	;
				tuser_save	[	124	]	<=	128'd0	;
				tuser_save	[	125	]	<=	128'd0	;
				tuser_save	[	126	]	<=	128'd0	;
				tuser_save	[	127	]	<=	128'd0	;
				tuser_save	[	128	]	<=	128'd0	;
				tuser_save	[	129	]	<=	128'd0	;
				tuser_save	[	130	]	<=	128'd0	;
				tuser_save	[	131	]	<=	128'd0	;
				tuser_save	[	132	]	<=	128'd0	;
				tuser_save	[	133	]	<=	128'd0	;
				tuser_save	[	134	]	<=	128'd0	;
				tuser_save	[	135	]	<=	128'd0	;
				tuser_save	[	136	]	<=	128'd0	;
				tuser_save	[	137	]	<=	128'd0	;
				tuser_save	[	138	]	<=	128'd0	;
				tuser_save	[	139	]	<=	128'd0	;
				tuser_save	[	140	]	<=	128'd0	;
				tuser_save	[	141	]	<=	128'd0	;
				tuser_save	[	142	]	<=	128'd0	;
				tuser_save	[	143	]	<=	128'd0	;
				tuser_save	[	144	]	<=	128'd0	;
				tuser_save	[	145	]	<=	128'd0	;
				tuser_save	[	146	]	<=	128'd0	;
				tuser_save	[	147	]	<=	128'd0	;
				tuser_save	[	148	]	<=	128'd0	;
				tuser_save	[	149	]	<=	128'd0	;
				tuser_save	[	150	]	<=	128'd0	;
				tuser_save	[	151	]	<=	128'd0	;
				tuser_save	[	152	]	<=	128'd0	;
				tuser_save	[	153	]	<=	128'd0	;
				tuser_save	[	154	]	<=	128'd0	;
				tuser_save	[	155	]	<=	128'd0	;
				tuser_save	[	156	]	<=	128'd0	;
				tuser_save	[	157	]	<=	128'd0	;
				tuser_save	[	158	]	<=	128'd0	;
				tuser_save	[	159	]	<=	128'd0	;
				tuser_save	[	160	]	<=	128'd0	;
				tuser_save	[	161	]	<=	128'd0	;
				tuser_save	[	162	]	<=	128'd0	;
				tuser_save	[	163	]	<=	128'd0	;
				tuser_save	[	164	]	<=	128'd0	;
				tuser_save	[	165	]	<=	128'd0	;
				tuser_save	[	166	]	<=	128'd0	;
				tuser_save	[	167	]	<=	128'd0	;
				tuser_save	[	168	]	<=	128'd0	;
				tuser_save	[	169	]	<=	128'd0	;
				tuser_save	[	170	]	<=	128'd0	;
				tuser_save	[	171	]	<=	128'd0	;
				tuser_save	[	172	]	<=	128'd0	;
				tuser_save	[	173	]	<=	128'd0	;
				tuser_save	[	174	]	<=	128'd0	;
				tuser_save	[	175	]	<=	128'd0	;
				tuser_save	[	176	]	<=	128'd0	;
				tuser_save	[	177	]	<=	128'd0	;
				tuser_save	[	178	]	<=	128'd0	;
				tuser_save	[	179	]	<=	128'd0	;
				tuser_save	[	180	]	<=	128'd0	;
				tuser_save	[	181	]	<=	128'd0	;
				tuser_save	[	182	]	<=	128'd0	;
				tuser_save	[	183	]	<=	128'd0	;
				tuser_save	[	184	]	<=	128'd0	;
				tuser_save	[	185	]	<=	128'd0	;
				tuser_save	[	186	]	<=	128'd0	;
				tuser_save	[	187	]	<=	128'd0	;
				tuser_save	[	188	]	<=	128'd0	;
				tuser_save	[	189	]	<=	128'd0	;
				tuser_save	[	190	]	<=	128'd0	;
				tuser_save	[	191	]	<=	128'd0	;
				tuser_save	[	192	]	<=	128'd0	;
				tuser_save	[	193	]	<=	128'd0	;
				tuser_save	[	194	]	<=	128'd0	;
				tuser_save	[	195	]	<=	128'd0	;
				tuser_save	[	196	]	<=	128'd0	;
				tuser_save	[	197	]	<=	128'd0	;
				tuser_save	[	198	]	<=	128'd0	;
				tuser_save	[	199	]	<=	128'd0	;
				tuser_save	[	200	]	<=	128'd0	;
				tuser_save	[	201	]	<=	128'd0	;
				tuser_save	[	202	]	<=	128'd0	;
				tuser_save	[	203	]	<=	128'd0	;
				tuser_save	[	204	]	<=	128'd0	;
				tuser_save	[	205	]	<=	128'd0	;
				tuser_save	[	206	]	<=	128'd0	;
				tuser_save	[	207	]	<=	128'd0	;
				tuser_save	[	208	]	<=	128'd0	;
				tuser_save	[	209	]	<=	128'd0	;
				tuser_save	[	210	]	<=	128'd0	;
				tuser_save	[	211	]	<=	128'd0	;
				tuser_save	[	212	]	<=	128'd0	;
				tuser_save	[	213	]	<=	128'd0	;
				tuser_save	[	214	]	<=	128'd0	;
				tuser_save	[	215	]	<=	128'd0	;
				tuser_save	[	216	]	<=	128'd0	;
				tuser_save	[	217	]	<=	128'd0	;
				tuser_save	[	218	]	<=	128'd0	;
				tuser_save	[	219	]	<=	128'd0	;
				tuser_save	[	220	]	<=	128'd0	;
				tuser_save	[	221	]	<=	128'd0	;
				tuser_save	[	222	]	<=	128'd0	;
				tuser_save	[	223	]	<=	128'd0	;
				tuser_save	[	224	]	<=	128'd0	;
				tuser_save	[	225	]	<=	128'd0	;
				tuser_save	[	226	]	<=	128'd0	;
				tuser_save	[	227	]	<=	128'd0	;
				tuser_save	[	228	]	<=	128'd0	;
				tuser_save	[	229	]	<=	128'd0	;
				tuser_save	[	230	]	<=	128'd0	;
				tuser_save	[	231	]	<=	128'd0	;
				tuser_save	[	232	]	<=	128'd0	;
				tuser_save	[	233	]	<=	128'd0	;
				tuser_save	[	234	]	<=	128'd0	;
				tuser_save	[	235	]	<=	128'd0	;
				tuser_save	[	236	]	<=	128'd0	;
				tuser_save	[	237	]	<=	128'd0	;
				tuser_save	[	238	]	<=	128'd0	;
				tuser_save	[	239	]	<=	128'd0	;
				tuser_save	[	240	]	<=	128'd0	;
				tuser_save	[	241	]	<=	128'd0	;
				tuser_save	[	242	]	<=	128'd0	;
				tuser_save	[	243	]	<=	128'd0	;
				tuser_save	[	244	]	<=	128'd0	;
				tuser_save	[	245	]	<=	128'd0	;
				tuser_save	[	246	]	<=	128'd0	;
				tuser_save	[	247	]	<=	128'd0	;
				tuser_save	[	248	]	<=	128'd0	;
				tuser_save	[	249	]	<=	128'd0	;
				tuser_save	[	250	]	<=	128'd0	;
				tuser_save	[	251	]	<=	128'd0	;
				tuser_save	[	252	]	<=	128'd0	;
				tuser_save	[	253	]	<=	128'd0	;
				tuser_save	[	254	]	<=	128'd0	;
				tuser_save	[	255	]	<=	128'd0	;
			count_packet	<= 2'd0;
			sum_tdata		<=	201'd0;
			sum_tuser		<=	128'd0;
			sum_tdata_valid		<=	1'b0;
			sum_tuser_valid		<=	1'b0;
			packet_num_count	<=	9'd0;
		end
		else if(axififo_din_valid)
		begin
			if(eth_type == 16'h0800)
			begin
				packet_num_count <= packet_num_count + 1'b1;
			end
			else
			begin
				packet_num_count <= packet_num_count;
			end
			if(tdata_save[255] == 201'd0)
			begin
				if((eth_type == 16'h0800) && (count_packet == 2'd0))
				begin
					tdata_save	[	0	]	<=	axififo_din;	//shift			
					tdata_save	[	1	]	<=	tdata_save	[	0	]	;
					tdata_save	[	2	]	<=	tdata_save	[	1	]	;
					tdata_save	[	3	]	<=	tdata_save	[	2	]	;
					tdata_save	[	4	]	<=	tdata_save	[	3	]	;
					tdata_save	[	5	]	<=	tdata_save	[	4	]	;
					tdata_save	[	6	]	<=	tdata_save	[	5	]	;
					tdata_save	[	7	]	<=	tdata_save	[	6	]	;
					tdata_save	[	8	]	<=	tdata_save	[	7	]	;
					tdata_save	[	9	]	<=	tdata_save	[	8	]	;
					tdata_save	[	10	]	<=	tdata_save	[	9	]	;
					tdata_save	[	11	]	<=	tdata_save	[	10	]	;
					tdata_save	[	12	]	<=	tdata_save	[	11	]	;
					tdata_save	[	13	]	<=	tdata_save	[	12	]	;
					tdata_save	[	14	]	<=	tdata_save	[	13	]	;
					tdata_save	[	15	]	<=	tdata_save	[	14	]	;
					tdata_save	[	16	]	<=	tdata_save	[	15	]	;
					tdata_save	[	17	]	<=	tdata_save	[	16	]	;
					tdata_save	[	18	]	<=	tdata_save	[	17	]	;
					tdata_save	[	19	]	<=	tdata_save	[	18	]	;
					tdata_save	[	20	]	<=	tdata_save	[	19	]	;
					tdata_save	[	21	]	<=	tdata_save	[	20	]	;
					tdata_save	[	22	]	<=	tdata_save	[	21	]	;
					tdata_save	[	23	]	<=	tdata_save	[	22	]	;
					tdata_save	[	24	]	<=	tdata_save	[	23	]	;
					tdata_save	[	25	]	<=	tdata_save	[	24	]	;
					tdata_save	[	26	]	<=	tdata_save	[	25	]	;
					tdata_save	[	27	]	<=	tdata_save	[	26	]	;
					tdata_save	[	28	]	<=	tdata_save	[	27	]	;
					tdata_save	[	29	]	<=	tdata_save	[	28	]	;
					tdata_save	[	30	]	<=	tdata_save	[	29	]	;
					tdata_save	[	31	]	<=	tdata_save	[	30	]	;
					tdata_save	[	32	]	<=	tdata_save	[	31	]	;
					tdata_save	[	33	]	<=	tdata_save	[	32	]	;
					tdata_save	[	34	]	<=	tdata_save	[	33	]	;
					tdata_save	[	35	]	<=	tdata_save	[	34	]	;
					tdata_save	[	36	]	<=	tdata_save	[	35	]	;
					tdata_save	[	37	]	<=	tdata_save	[	36	]	;
					tdata_save	[	38	]	<=	tdata_save	[	37	]	;
					tdata_save	[	39	]	<=	tdata_save	[	38	]	;
					tdata_save	[	40	]	<=	tdata_save	[	39	]	;
					tdata_save	[	41	]	<=	tdata_save	[	40	]	;
					tdata_save	[	42	]	<=	tdata_save	[	41	]	;
					tdata_save	[	43	]	<=	tdata_save	[	42	]	;
					tdata_save	[	44	]	<=	tdata_save	[	43	]	;
					tdata_save	[	45	]	<=	tdata_save	[	44	]	;
					tdata_save	[	46	]	<=	tdata_save	[	45	]	;
					tdata_save	[	47	]	<=	tdata_save	[	46	]	;
					tdata_save	[	48	]	<=	tdata_save	[	47	]	;
					tdata_save	[	49	]	<=	tdata_save	[	48	]	;
					tdata_save	[	50	]	<=	tdata_save	[	49	]	;
					tdata_save	[	51	]	<=	tdata_save	[	50	]	;
					tdata_save	[	52	]	<=	tdata_save	[	51	]	;
					tdata_save	[	53	]	<=	tdata_save	[	52	]	;
					tdata_save	[	54	]	<=	tdata_save	[	53	]	;
					tdata_save	[	55	]	<=	tdata_save	[	54	]	;
					tdata_save	[	56	]	<=	tdata_save	[	55	]	;
					tdata_save	[	57	]	<=	tdata_save	[	56	]	;
					tdata_save	[	58	]	<=	tdata_save	[	57	]	;
					tdata_save	[	59	]	<=	tdata_save	[	58	]	;
					tdata_save	[	60	]	<=	tdata_save	[	59	]	;
					tdata_save	[	61	]	<=	tdata_save	[	60	]	;
					tdata_save	[	62	]	<=	tdata_save	[	61	]	;
					tdata_save	[	63	]	<=	tdata_save	[	62	]	;
					tdata_save	[	64	]	<=	tdata_save	[	63	]	;
					tdata_save	[	65	]	<=	tdata_save	[	64	]	;
					tdata_save	[	66	]	<=	tdata_save	[	65	]	;
					tdata_save	[	67	]	<=	tdata_save	[	66	]	;
					tdata_save	[	68	]	<=	tdata_save	[	67	]	;
					tdata_save	[	69	]	<=	tdata_save	[	68	]	;
					tdata_save	[	70	]	<=	tdata_save	[	69	]	;
					tdata_save	[	71	]	<=	tdata_save	[	70	]	;
					tdata_save	[	72	]	<=	tdata_save	[	71	]	;
					tdata_save	[	73	]	<=	tdata_save	[	72	]	;
					tdata_save	[	74	]	<=	tdata_save	[	73	]	;
					tdata_save	[	75	]	<=	tdata_save	[	74	]	;
					tdata_save	[	76	]	<=	tdata_save	[	75	]	;
					tdata_save	[	77	]	<=	tdata_save	[	76	]	;
					tdata_save	[	78	]	<=	tdata_save	[	77	]	;
					tdata_save	[	79	]	<=	tdata_save	[	78	]	;
					tdata_save	[	80	]	<=	tdata_save	[	79	]	;
					tdata_save	[	81	]	<=	tdata_save	[	80	]	;
					tdata_save	[	82	]	<=	tdata_save	[	81	]	;
					tdata_save	[	83	]	<=	tdata_save	[	82	]	;
					tdata_save	[	84	]	<=	tdata_save	[	83	]	;
					tdata_save	[	85	]	<=	tdata_save	[	84	]	;
					tdata_save	[	86	]	<=	tdata_save	[	85	]	;
					tdata_save	[	87	]	<=	tdata_save	[	86	]	;
					tdata_save	[	88	]	<=	tdata_save	[	87	]	;
					tdata_save	[	89	]	<=	tdata_save	[	88	]	;
					tdata_save	[	90	]	<=	tdata_save	[	89	]	;
					tdata_save	[	91	]	<=	tdata_save	[	90	]	;
					tdata_save	[	92	]	<=	tdata_save	[	91	]	;
					tdata_save	[	93	]	<=	tdata_save	[	92	]	;
					tdata_save	[	94	]	<=	tdata_save	[	93	]	;
					tdata_save	[	95	]	<=	tdata_save	[	94	]	;
					tdata_save	[	96	]	<=	tdata_save	[	95	]	;
					tdata_save	[	97	]	<=	tdata_save	[	96	]	;
					tdata_save	[	98	]	<=	tdata_save	[	97	]	;
					tdata_save	[	99	]	<=	tdata_save	[	98	]	;
					tdata_save	[	100	]	<=	tdata_save	[	99	]	;
					tdata_save	[	101	]	<=	tdata_save	[	100	]	;
					tdata_save	[	102	]	<=	tdata_save	[	101	]	;
					tdata_save	[	103	]	<=	tdata_save	[	102	]	;
					tdata_save	[	104	]	<=	tdata_save	[	103	]	;
					tdata_save	[	105	]	<=	tdata_save	[	104	]	;
					tdata_save	[	106	]	<=	tdata_save	[	105	]	;
					tdata_save	[	107	]	<=	tdata_save	[	106	]	;
					tdata_save	[	108	]	<=	tdata_save	[	107	]	;
					tdata_save	[	109	]	<=	tdata_save	[	108	]	;
					tdata_save	[	110	]	<=	tdata_save	[	109	]	;
					tdata_save	[	111	]	<=	tdata_save	[	110	]	;
					tdata_save	[	112	]	<=	tdata_save	[	111	]	;
					tdata_save	[	113	]	<=	tdata_save	[	112	]	;
					tdata_save	[	114	]	<=	tdata_save	[	113	]	;
					tdata_save	[	115	]	<=	tdata_save	[	114	]	;
					tdata_save	[	116	]	<=	tdata_save	[	115	]	;
					tdata_save	[	117	]	<=	tdata_save	[	116	]	;
					tdata_save	[	118	]	<=	tdata_save	[	117	]	;
					tdata_save	[	119	]	<=	tdata_save	[	118	]	;
					tdata_save	[	120	]	<=	tdata_save	[	119	]	;
					tdata_save	[	121	]	<=	tdata_save	[	120	]	;
					tdata_save	[	122	]	<=	tdata_save	[	121	]	;
					tdata_save	[	123	]	<=	tdata_save	[	122	]	;
					tdata_save	[	124	]	<=	tdata_save	[	123	]	;
					tdata_save	[	125	]	<=	tdata_save	[	124	]	;
					tdata_save	[	126	]	<=	tdata_save	[	125	]	;
					tdata_save	[	127	]	<=	tdata_save	[	126	]	;
					tdata_save	[	128	]	<=	tdata_save	[	127	]	;
					tdata_save	[	129	]	<=	tdata_save	[	128	]	;
					tdata_save	[	130	]	<=	tdata_save	[	129	]	;
					tdata_save	[	131	]	<=	tdata_save	[	130	]	;
					tdata_save	[	132	]	<=	tdata_save	[	131	]	;
					tdata_save	[	133	]	<=	tdata_save	[	132	]	;
					tdata_save	[	134	]	<=	tdata_save	[	133	]	;
					tdata_save	[	135	]	<=	tdata_save	[	134	]	;
					tdata_save	[	136	]	<=	tdata_save	[	135	]	;
					tdata_save	[	137	]	<=	tdata_save	[	136	]	;
					tdata_save	[	138	]	<=	tdata_save	[	137	]	;
					tdata_save	[	139	]	<=	tdata_save	[	138	]	;
					tdata_save	[	140	]	<=	tdata_save	[	139	]	;
					tdata_save	[	141	]	<=	tdata_save	[	140	]	;
					tdata_save	[	142	]	<=	tdata_save	[	141	]	;
					tdata_save	[	143	]	<=	tdata_save	[	142	]	;
					tdata_save	[	144	]	<=	tdata_save	[	143	]	;
					tdata_save	[	145	]	<=	tdata_save	[	144	]	;
					tdata_save	[	146	]	<=	tdata_save	[	145	]	;
					tdata_save	[	147	]	<=	tdata_save	[	146	]	;
					tdata_save	[	148	]	<=	tdata_save	[	147	]	;
					tdata_save	[	149	]	<=	tdata_save	[	148	]	;
					tdata_save	[	150	]	<=	tdata_save	[	149	]	;
					tdata_save	[	151	]	<=	tdata_save	[	150	]	;
					tdata_save	[	152	]	<=	tdata_save	[	151	]	;
					tdata_save	[	153	]	<=	tdata_save	[	152	]	;
					tdata_save	[	154	]	<=	tdata_save	[	153	]	;
					tdata_save	[	155	]	<=	tdata_save	[	154	]	;
					tdata_save	[	156	]	<=	tdata_save	[	155	]	;
					tdata_save	[	157	]	<=	tdata_save	[	156	]	;
					tdata_save	[	158	]	<=	tdata_save	[	157	]	;
					tdata_save	[	159	]	<=	tdata_save	[	158	]	;
					tdata_save	[	160	]	<=	tdata_save	[	159	]	;
					tdata_save	[	161	]	<=	tdata_save	[	160	]	;
					tdata_save	[	162	]	<=	tdata_save	[	161	]	;
					tdata_save	[	163	]	<=	tdata_save	[	162	]	;
					tdata_save	[	164	]	<=	tdata_save	[	163	]	;
					tdata_save	[	165	]	<=	tdata_save	[	164	]	;
					tdata_save	[	166	]	<=	tdata_save	[	165	]	;
					tdata_save	[	167	]	<=	tdata_save	[	166	]	;
					tdata_save	[	168	]	<=	tdata_save	[	167	]	;
					tdata_save	[	169	]	<=	tdata_save	[	168	]	;
					tdata_save	[	170	]	<=	tdata_save	[	169	]	;
					tdata_save	[	171	]	<=	tdata_save	[	170	]	;
					tdata_save	[	172	]	<=	tdata_save	[	171	]	;
					tdata_save	[	173	]	<=	tdata_save	[	172	]	;
					tdata_save	[	174	]	<=	tdata_save	[	173	]	;
					tdata_save	[	175	]	<=	tdata_save	[	174	]	;
					tdata_save	[	176	]	<=	tdata_save	[	175	]	;
					tdata_save	[	177	]	<=	tdata_save	[	176	]	;
					tdata_save	[	178	]	<=	tdata_save	[	177	]	;
					tdata_save	[	179	]	<=	tdata_save	[	178	]	;
					tdata_save	[	180	]	<=	tdata_save	[	179	]	;
					tdata_save	[	181	]	<=	tdata_save	[	180	]	;
					tdata_save	[	182	]	<=	tdata_save	[	181	]	;
					tdata_save	[	183	]	<=	tdata_save	[	182	]	;
					tdata_save	[	184	]	<=	tdata_save	[	183	]	;
					tdata_save	[	185	]	<=	tdata_save	[	184	]	;
					tdata_save	[	186	]	<=	tdata_save	[	185	]	;
					tdata_save	[	187	]	<=	tdata_save	[	186	]	;
					tdata_save	[	188	]	<=	tdata_save	[	187	]	;
					tdata_save	[	189	]	<=	tdata_save	[	188	]	;
					tdata_save	[	190	]	<=	tdata_save	[	189	]	;
					tdata_save	[	191	]	<=	tdata_save	[	190	]	;
					tdata_save	[	192	]	<=	tdata_save	[	191	]	;
					tdata_save	[	193	]	<=	tdata_save	[	192	]	;
					tdata_save	[	194	]	<=	tdata_save	[	193	]	;
					tdata_save	[	195	]	<=	tdata_save	[	194	]	;
					tdata_save	[	196	]	<=	tdata_save	[	195	]	;
					tdata_save	[	197	]	<=	tdata_save	[	196	]	;
					tdata_save	[	198	]	<=	tdata_save	[	197	]	;
					tdata_save	[	199	]	<=	tdata_save	[	198	]	;
					tdata_save	[	200	]	<=	tdata_save	[	199	]	;
					tdata_save	[	201	]	<=	tdata_save	[	200	]	;
					tdata_save	[	202	]	<=	tdata_save	[	201	]	;
					tdata_save	[	203	]	<=	tdata_save	[	202	]	;
					tdata_save	[	204	]	<=	tdata_save	[	203	]	;
					tdata_save	[	205	]	<=	tdata_save	[	204	]	;
					tdata_save	[	206	]	<=	tdata_save	[	205	]	;
					tdata_save	[	207	]	<=	tdata_save	[	206	]	;
					tdata_save	[	208	]	<=	tdata_save	[	207	]	;
					tdata_save	[	209	]	<=	tdata_save	[	208	]	;
					tdata_save	[	210	]	<=	tdata_save	[	209	]	;
					tdata_save	[	211	]	<=	tdata_save	[	210	]	;
					tdata_save	[	212	]	<=	tdata_save	[	211	]	;
					tdata_save	[	213	]	<=	tdata_save	[	212	]	;
					tdata_save	[	214	]	<=	tdata_save	[	213	]	;
					tdata_save	[	215	]	<=	tdata_save	[	214	]	;
					tdata_save	[	216	]	<=	tdata_save	[	215	]	;
					tdata_save	[	217	]	<=	tdata_save	[	216	]	;
					tdata_save	[	218	]	<=	tdata_save	[	217	]	;
					tdata_save	[	219	]	<=	tdata_save	[	218	]	;
					tdata_save	[	220	]	<=	tdata_save	[	219	]	;
					tdata_save	[	221	]	<=	tdata_save	[	220	]	;
					tdata_save	[	222	]	<=	tdata_save	[	221	]	;
					tdata_save	[	223	]	<=	tdata_save	[	222	]	;
					tdata_save	[	224	]	<=	tdata_save	[	223	]	;
					tdata_save	[	225	]	<=	tdata_save	[	224	]	;
					tdata_save	[	226	]	<=	tdata_save	[	225	]	;
					tdata_save	[	227	]	<=	tdata_save	[	226	]	;
					tdata_save	[	228	]	<=	tdata_save	[	227	]	;
					tdata_save	[	229	]	<=	tdata_save	[	228	]	;
					tdata_save	[	230	]	<=	tdata_save	[	229	]	;
					tdata_save	[	231	]	<=	tdata_save	[	230	]	;
					tdata_save	[	232	]	<=	tdata_save	[	231	]	;
					tdata_save	[	233	]	<=	tdata_save	[	232	]	;
					tdata_save	[	234	]	<=	tdata_save	[	233	]	;
					tdata_save	[	235	]	<=	tdata_save	[	234	]	;
					tdata_save	[	236	]	<=	tdata_save	[	235	]	;
					tdata_save	[	237	]	<=	tdata_save	[	236	]	;
					tdata_save	[	238	]	<=	tdata_save	[	237	]	;
					tdata_save	[	239	]	<=	tdata_save	[	238	]	;
					tdata_save	[	240	]	<=	tdata_save	[	239	]	;
					tdata_save	[	241	]	<=	tdata_save	[	240	]	;
					tdata_save	[	242	]	<=	tdata_save	[	241	]	;
					tdata_save	[	243	]	<=	tdata_save	[	242	]	;
					tdata_save	[	244	]	<=	tdata_save	[	243	]	;
					tdata_save	[	245	]	<=	tdata_save	[	244	]	;
					tdata_save	[	246	]	<=	tdata_save	[	245	]	;
					tdata_save	[	247	]	<=	tdata_save	[	246	]	;
					tdata_save	[	248	]	<=	tdata_save	[	247	]	;
					tdata_save	[	249	]	<=	tdata_save	[	248	]	;
					tdata_save	[	250	]	<=	tdata_save	[	249	]	;
					tdata_save	[	251	]	<=	tdata_save	[	250	]	;
					tdata_save	[	252	]	<=	tdata_save	[	251	]	;
					tdata_save	[	253	]	<=	tdata_save	[	252	]	;
					tdata_save	[	254	]	<=	tdata_save	[	253	]	;
					tdata_save	[	255	]	<=	tdata_save	[	254	]	;
					tuser_save	[	0	]	<=	tuser;						
				tuser_save	[	1	]	<=	tuser_save	[	0	]	;
				tuser_save	[	2	]	<=	tuser_save	[	1	]	;
				tuser_save	[	3	]	<=	tuser_save	[	2	]	;
				tuser_save	[	4	]	<=	tuser_save	[	3	]	;
				tuser_save	[	5	]	<=	tuser_save	[	4	]	;
				tuser_save	[	6	]	<=	tuser_save	[	5	]	;
				tuser_save	[	7	]	<=	tuser_save	[	6	]	;
				tuser_save	[	8	]	<=	tuser_save	[	7	]	;
				tuser_save	[	9	]	<=	tuser_save	[	8	]	;
				tuser_save	[	10	]	<=	tuser_save	[	9	]	;
				tuser_save	[	11	]	<=	tuser_save	[	10	]	;
				tuser_save	[	12	]	<=	tuser_save	[	11	]	;
				tuser_save	[	13	]	<=	tuser_save	[	12	]	;
				tuser_save	[	14	]	<=	tuser_save	[	13	]	;
				tuser_save	[	15	]	<=	tuser_save	[	14	]	;
				tuser_save	[	16	]	<=	tuser_save	[	15	]	;
				tuser_save	[	17	]	<=	tuser_save	[	16	]	;
				tuser_save	[	18	]	<=	tuser_save	[	17	]	;
				tuser_save	[	19	]	<=	tuser_save	[	18	]	;
				tuser_save	[	20	]	<=	tuser_save	[	19	]	;
				tuser_save	[	21	]	<=	tuser_save	[	20	]	;
				tuser_save	[	22	]	<=	tuser_save	[	21	]	;
				tuser_save	[	23	]	<=	tuser_save	[	22	]	;
				tuser_save	[	24	]	<=	tuser_save	[	23	]	;
				tuser_save	[	25	]	<=	tuser_save	[	24	]	;
				tuser_save	[	26	]	<=	tuser_save	[	25	]	;
				tuser_save	[	27	]	<=	tuser_save	[	26	]	;
				tuser_save	[	28	]	<=	tuser_save	[	27	]	;
				tuser_save	[	29	]	<=	tuser_save	[	28	]	;
				tuser_save	[	30	]	<=	tuser_save	[	29	]	;
				tuser_save	[	31	]	<=	tuser_save	[	30	]	;
				tuser_save	[	32	]	<=	tuser_save	[	31	]	;
				tuser_save	[	33	]	<=	tuser_save	[	32	]	;
				tuser_save	[	34	]	<=	tuser_save	[	33	]	;
				tuser_save	[	35	]	<=	tuser_save	[	34	]	;
				tuser_save	[	36	]	<=	tuser_save	[	35	]	;
				tuser_save	[	37	]	<=	tuser_save	[	36	]	;
				tuser_save	[	38	]	<=	tuser_save	[	37	]	;
				tuser_save	[	39	]	<=	tuser_save	[	38	]	;
				tuser_save	[	40	]	<=	tuser_save	[	39	]	;
				tuser_save	[	41	]	<=	tuser_save	[	40	]	;
				tuser_save	[	42	]	<=	tuser_save	[	41	]	;
				tuser_save	[	43	]	<=	tuser_save	[	42	]	;
				tuser_save	[	44	]	<=	tuser_save	[	43	]	;
				tuser_save	[	45	]	<=	tuser_save	[	44	]	;
				tuser_save	[	46	]	<=	tuser_save	[	45	]	;
				tuser_save	[	47	]	<=	tuser_save	[	46	]	;
				tuser_save	[	48	]	<=	tuser_save	[	47	]	;
				tuser_save	[	49	]	<=	tuser_save	[	48	]	;
				tuser_save	[	50	]	<=	tuser_save	[	49	]	;
				tuser_save	[	51	]	<=	tuser_save	[	50	]	;
				tuser_save	[	52	]	<=	tuser_save	[	51	]	;
				tuser_save	[	53	]	<=	tuser_save	[	52	]	;
				tuser_save	[	54	]	<=	tuser_save	[	53	]	;
				tuser_save	[	55	]	<=	tuser_save	[	54	]	;
				tuser_save	[	56	]	<=	tuser_save	[	55	]	;
				tuser_save	[	57	]	<=	tuser_save	[	56	]	;
				tuser_save	[	58	]	<=	tuser_save	[	57	]	;
				tuser_save	[	59	]	<=	tuser_save	[	58	]	;
				tuser_save	[	60	]	<=	tuser_save	[	59	]	;
				tuser_save	[	61	]	<=	tuser_save	[	60	]	;
				tuser_save	[	62	]	<=	tuser_save	[	61	]	;
				tuser_save	[	63	]	<=	tuser_save	[	62	]	;
				tuser_save	[	64	]	<=	tuser_save	[	63	]	;
				tuser_save	[	65	]	<=	tuser_save	[	64	]	;
				tuser_save	[	66	]	<=	tuser_save	[	65	]	;
				tuser_save	[	67	]	<=	tuser_save	[	66	]	;
				tuser_save	[	68	]	<=	tuser_save	[	67	]	;
				tuser_save	[	69	]	<=	tuser_save	[	68	]	;
				tuser_save	[	70	]	<=	tuser_save	[	69	]	;
				tuser_save	[	71	]	<=	tuser_save	[	70	]	;
				tuser_save	[	72	]	<=	tuser_save	[	71	]	;
				tuser_save	[	73	]	<=	tuser_save	[	72	]	;
				tuser_save	[	74	]	<=	tuser_save	[	73	]	;
				tuser_save	[	75	]	<=	tuser_save	[	74	]	;
				tuser_save	[	76	]	<=	tuser_save	[	75	]	;
				tuser_save	[	77	]	<=	tuser_save	[	76	]	;
				tuser_save	[	78	]	<=	tuser_save	[	77	]	;
				tuser_save	[	79	]	<=	tuser_save	[	78	]	;
				tuser_save	[	80	]	<=	tuser_save	[	79	]	;
				tuser_save	[	81	]	<=	tuser_save	[	80	]	;
				tuser_save	[	82	]	<=	tuser_save	[	81	]	;
				tuser_save	[	83	]	<=	tuser_save	[	82	]	;
				tuser_save	[	84	]	<=	tuser_save	[	83	]	;
				tuser_save	[	85	]	<=	tuser_save	[	84	]	;
				tuser_save	[	86	]	<=	tuser_save	[	85	]	;
				tuser_save	[	87	]	<=	tuser_save	[	86	]	;
				tuser_save	[	88	]	<=	tuser_save	[	87	]	;
				tuser_save	[	89	]	<=	tuser_save	[	88	]	;
				tuser_save	[	90	]	<=	tuser_save	[	89	]	;
				tuser_save	[	91	]	<=	tuser_save	[	90	]	;
				tuser_save	[	92	]	<=	tuser_save	[	91	]	;
				tuser_save	[	93	]	<=	tuser_save	[	92	]	;
				tuser_save	[	94	]	<=	tuser_save	[	93	]	;
				tuser_save	[	95	]	<=	tuser_save	[	94	]	;
				tuser_save	[	96	]	<=	tuser_save	[	95	]	;
				tuser_save	[	97	]	<=	tuser_save	[	96	]	;
				tuser_save	[	98	]	<=	tuser_save	[	97	]	;
				tuser_save	[	99	]	<=	tuser_save	[	98	]	;
				tuser_save	[	100	]	<=	tuser_save	[	99	]	;
				tuser_save	[	101	]	<=	tuser_save	[	100	]	;
				tuser_save	[	102	]	<=	tuser_save	[	101	]	;
				tuser_save	[	103	]	<=	tuser_save	[	102	]	;
				tuser_save	[	104	]	<=	tuser_save	[	103	]	;
				tuser_save	[	105	]	<=	tuser_save	[	104	]	;
				tuser_save	[	106	]	<=	tuser_save	[	105	]	;
				tuser_save	[	107	]	<=	tuser_save	[	106	]	;
				tuser_save	[	108	]	<=	tuser_save	[	107	]	;
				tuser_save	[	109	]	<=	tuser_save	[	108	]	;
				tuser_save	[	110	]	<=	tuser_save	[	109	]	;
				tuser_save	[	111	]	<=	tuser_save	[	110	]	;
				tuser_save	[	112	]	<=	tuser_save	[	111	]	;
				tuser_save	[	113	]	<=	tuser_save	[	112	]	;
				tuser_save	[	114	]	<=	tuser_save	[	113	]	;
				tuser_save	[	115	]	<=	tuser_save	[	114	]	;
				tuser_save	[	116	]	<=	tuser_save	[	115	]	;
				tuser_save	[	117	]	<=	tuser_save	[	116	]	;
				tuser_save	[	118	]	<=	tuser_save	[	117	]	;
				tuser_save	[	119	]	<=	tuser_save	[	118	]	;
				tuser_save	[	120	]	<=	tuser_save	[	119	]	;
				tuser_save	[	121	]	<=	tuser_save	[	120	]	;
				tuser_save	[	122	]	<=	tuser_save	[	121	]	;
				tuser_save	[	123	]	<=	tuser_save	[	122	]	;
				tuser_save	[	124	]	<=	tuser_save	[	123	]	;
				tuser_save	[	125	]	<=	tuser_save	[	124	]	;
				tuser_save	[	126	]	<=	tuser_save	[	125	]	;
				tuser_save	[	127	]	<=	tuser_save	[	126	]	;
				tuser_save	[	128	]	<=	tuser_save	[	127	]	;
				tuser_save	[	129	]	<=	tuser_save	[	128	]	;
				tuser_save	[	130	]	<=	tuser_save	[	129	]	;
				tuser_save	[	131	]	<=	tuser_save	[	130	]	;
				tuser_save	[	132	]	<=	tuser_save	[	131	]	;
				tuser_save	[	133	]	<=	tuser_save	[	132	]	;
				tuser_save	[	134	]	<=	tuser_save	[	133	]	;
				tuser_save	[	135	]	<=	tuser_save	[	134	]	;
				tuser_save	[	136	]	<=	tuser_save	[	135	]	;
				tuser_save	[	137	]	<=	tuser_save	[	136	]	;
				tuser_save	[	138	]	<=	tuser_save	[	137	]	;
				tuser_save	[	139	]	<=	tuser_save	[	138	]	;
				tuser_save	[	140	]	<=	tuser_save	[	139	]	;
				tuser_save	[	141	]	<=	tuser_save	[	140	]	;
				tuser_save	[	142	]	<=	tuser_save	[	141	]	;
				tuser_save	[	143	]	<=	tuser_save	[	142	]	;
				tuser_save	[	144	]	<=	tuser_save	[	143	]	;
				tuser_save	[	145	]	<=	tuser_save	[	144	]	;
				tuser_save	[	146	]	<=	tuser_save	[	145	]	;
				tuser_save	[	147	]	<=	tuser_save	[	146	]	;
				tuser_save	[	148	]	<=	tuser_save	[	147	]	;
				tuser_save	[	149	]	<=	tuser_save	[	148	]	;
				tuser_save	[	150	]	<=	tuser_save	[	149	]	;
				tuser_save	[	151	]	<=	tuser_save	[	150	]	;
				tuser_save	[	152	]	<=	tuser_save	[	151	]	;
				tuser_save	[	153	]	<=	tuser_save	[	152	]	;
				tuser_save	[	154	]	<=	tuser_save	[	153	]	;
				tuser_save	[	155	]	<=	tuser_save	[	154	]	;
				tuser_save	[	156	]	<=	tuser_save	[	155	]	;
				tuser_save	[	157	]	<=	tuser_save	[	156	]	;
				tuser_save	[	158	]	<=	tuser_save	[	157	]	;
				tuser_save	[	159	]	<=	tuser_save	[	158	]	;
				tuser_save	[	160	]	<=	tuser_save	[	159	]	;
				tuser_save	[	161	]	<=	tuser_save	[	160	]	;
				tuser_save	[	162	]	<=	tuser_save	[	161	]	;
				tuser_save	[	163	]	<=	tuser_save	[	162	]	;
				tuser_save	[	164	]	<=	tuser_save	[	163	]	;
				tuser_save	[	165	]	<=	tuser_save	[	164	]	;
				tuser_save	[	166	]	<=	tuser_save	[	165	]	;
				tuser_save	[	167	]	<=	tuser_save	[	166	]	;
				tuser_save	[	168	]	<=	tuser_save	[	167	]	;
				tuser_save	[	169	]	<=	tuser_save	[	168	]	;
				tuser_save	[	170	]	<=	tuser_save	[	169	]	;
				tuser_save	[	171	]	<=	tuser_save	[	170	]	;
				tuser_save	[	172	]	<=	tuser_save	[	171	]	;
				tuser_save	[	173	]	<=	tuser_save	[	172	]	;
				tuser_save	[	174	]	<=	tuser_save	[	173	]	;
				tuser_save	[	175	]	<=	tuser_save	[	174	]	;
				tuser_save	[	176	]	<=	tuser_save	[	175	]	;
				tuser_save	[	177	]	<=	tuser_save	[	176	]	;
				tuser_save	[	178	]	<=	tuser_save	[	177	]	;
				tuser_save	[	179	]	<=	tuser_save	[	178	]	;
				tuser_save	[	180	]	<=	tuser_save	[	179	]	;
				tuser_save	[	181	]	<=	tuser_save	[	180	]	;
				tuser_save	[	182	]	<=	tuser_save	[	181	]	;
				tuser_save	[	183	]	<=	tuser_save	[	182	]	;
				tuser_save	[	184	]	<=	tuser_save	[	183	]	;
				tuser_save	[	185	]	<=	tuser_save	[	184	]	;
				tuser_save	[	186	]	<=	tuser_save	[	185	]	;
				tuser_save	[	187	]	<=	tuser_save	[	186	]	;
				tuser_save	[	188	]	<=	tuser_save	[	187	]	;
				tuser_save	[	189	]	<=	tuser_save	[	188	]	;
				tuser_save	[	190	]	<=	tuser_save	[	189	]	;
				tuser_save	[	191	]	<=	tuser_save	[	190	]	;
				tuser_save	[	192	]	<=	tuser_save	[	191	]	;
				tuser_save	[	193	]	<=	tuser_save	[	192	]	;
				tuser_save	[	194	]	<=	tuser_save	[	193	]	;
				tuser_save	[	195	]	<=	tuser_save	[	194	]	;
				tuser_save	[	196	]	<=	tuser_save	[	195	]	;
				tuser_save	[	197	]	<=	tuser_save	[	196	]	;
				tuser_save	[	198	]	<=	tuser_save	[	197	]	;
				tuser_save	[	199	]	<=	tuser_save	[	198	]	;
				tuser_save	[	200	]	<=	tuser_save	[	199	]	;
				tuser_save	[	201	]	<=	tuser_save	[	200	]	;
				tuser_save	[	202	]	<=	tuser_save	[	201	]	;
				tuser_save	[	203	]	<=	tuser_save	[	202	]	;
				tuser_save	[	204	]	<=	tuser_save	[	203	]	;
				tuser_save	[	205	]	<=	tuser_save	[	204	]	;
				tuser_save	[	206	]	<=	tuser_save	[	205	]	;
				tuser_save	[	207	]	<=	tuser_save	[	206	]	;
				tuser_save	[	208	]	<=	tuser_save	[	207	]	;
				tuser_save	[	209	]	<=	tuser_save	[	208	]	;
				tuser_save	[	210	]	<=	tuser_save	[	209	]	;
				tuser_save	[	211	]	<=	tuser_save	[	210	]	;
				tuser_save	[	212	]	<=	tuser_save	[	211	]	;
				tuser_save	[	213	]	<=	tuser_save	[	212	]	;
				tuser_save	[	214	]	<=	tuser_save	[	213	]	;
				tuser_save	[	215	]	<=	tuser_save	[	214	]	;
				tuser_save	[	216	]	<=	tuser_save	[	215	]	;
				tuser_save	[	217	]	<=	tuser_save	[	216	]	;
				tuser_save	[	218	]	<=	tuser_save	[	217	]	;
				tuser_save	[	219	]	<=	tuser_save	[	218	]	;
				tuser_save	[	220	]	<=	tuser_save	[	219	]	;
				tuser_save	[	221	]	<=	tuser_save	[	220	]	;
				tuser_save	[	222	]	<=	tuser_save	[	221	]	;
				tuser_save	[	223	]	<=	tuser_save	[	222	]	;
				tuser_save	[	224	]	<=	tuser_save	[	223	]	;
				tuser_save	[	225	]	<=	tuser_save	[	224	]	;
				tuser_save	[	226	]	<=	tuser_save	[	225	]	;
				tuser_save	[	227	]	<=	tuser_save	[	226	]	;
				tuser_save	[	228	]	<=	tuser_save	[	227	]	;
				tuser_save	[	229	]	<=	tuser_save	[	228	]	;
				tuser_save	[	230	]	<=	tuser_save	[	229	]	;
				tuser_save	[	231	]	<=	tuser_save	[	230	]	;
				tuser_save	[	232	]	<=	tuser_save	[	231	]	;
				tuser_save	[	233	]	<=	tuser_save	[	232	]	;
				tuser_save	[	234	]	<=	tuser_save	[	233	]	;
				tuser_save	[	235	]	<=	tuser_save	[	234	]	;
				tuser_save	[	236	]	<=	tuser_save	[	235	]	;
				tuser_save	[	237	]	<=	tuser_save	[	236	]	;
				tuser_save	[	238	]	<=	tuser_save	[	237	]	;
				tuser_save	[	239	]	<=	tuser_save	[	238	]	;
				tuser_save	[	240	]	<=	tuser_save	[	239	]	;
				tuser_save	[	241	]	<=	tuser_save	[	240	]	;
				tuser_save	[	242	]	<=	tuser_save	[	241	]	;
				tuser_save	[	243	]	<=	tuser_save	[	242	]	;
				tuser_save	[	244	]	<=	tuser_save	[	243	]	;
				tuser_save	[	245	]	<=	tuser_save	[	244	]	;
				tuser_save	[	246	]	<=	tuser_save	[	245	]	;
				tuser_save	[	247	]	<=	tuser_save	[	246	]	;
				tuser_save	[	248	]	<=	tuser_save	[	247	]	;
				tuser_save	[	249	]	<=	tuser_save	[	248	]	;
				tuser_save	[	250	]	<=	tuser_save	[	249	]	;
				tuser_save	[	251	]	<=	tuser_save	[	250	]	;
				tuser_save	[	252	]	<=	tuser_save	[	251	]	;
				tuser_save	[	253	]	<=	tuser_save	[	252	]	;
				tuser_save	[	254	]	<=	tuser_save	[	253	]	;
				tuser_save	[	255	]	<=	tuser_save	[	254	]	;
					if(count_packet == 2'd2)
					begin
						count_packet <= 2'd0;
					end
					else
					begin
						count_packet	<= count_packet + 1'b1;
					end
					sum_tdata		<=	201'd0;
					sum_tuser		<=	128'd0;
					sum_tdata_valid		<=	1'b0;
					sum_tuser_valid		<=	1'b0;
				end
				else if(count_packet == 2'd1)
				begin
					tdata_save	[	0	]	<=	axififo_din;	//shift			
					tdata_save	[	1	]	<=	tdata_save	[	0	]	;
					tdata_save	[	2	]	<=	tdata_save	[	1	]	;
					tdata_save	[	3	]	<=	tdata_save	[	2	]	;
					tdata_save	[	4	]	<=	tdata_save	[	3	]	;
					tdata_save	[	5	]	<=	tdata_save	[	4	]	;
					tdata_save	[	6	]	<=	tdata_save	[	5	]	;
					tdata_save	[	7	]	<=	tdata_save	[	6	]	;
					tdata_save	[	8	]	<=	tdata_save	[	7	]	;
					tdata_save	[	9	]	<=	tdata_save	[	8	]	;
					tdata_save	[	10	]	<=	tdata_save	[	9	]	;
					tdata_save	[	11	]	<=	tdata_save	[	10	]	;
					tdata_save	[	12	]	<=	tdata_save	[	11	]	;
					tdata_save	[	13	]	<=	tdata_save	[	12	]	;
					tdata_save	[	14	]	<=	tdata_save	[	13	]	;
					tdata_save	[	15	]	<=	tdata_save	[	14	]	;
					tdata_save	[	16	]	<=	tdata_save	[	15	]	;
					tdata_save	[	17	]	<=	tdata_save	[	16	]	;
					tdata_save	[	18	]	<=	tdata_save	[	17	]	;
					tdata_save	[	19	]	<=	tdata_save	[	18	]	;
					tdata_save	[	20	]	<=	tdata_save	[	19	]	;
					tdata_save	[	21	]	<=	tdata_save	[	20	]	;
					tdata_save	[	22	]	<=	tdata_save	[	21	]	;
					tdata_save	[	23	]	<=	tdata_save	[	22	]	;
					tdata_save	[	24	]	<=	tdata_save	[	23	]	;
					tdata_save	[	25	]	<=	tdata_save	[	24	]	;
					tdata_save	[	26	]	<=	tdata_save	[	25	]	;
					tdata_save	[	27	]	<=	tdata_save	[	26	]	;
					tdata_save	[	28	]	<=	tdata_save	[	27	]	;
					tdata_save	[	29	]	<=	tdata_save	[	28	]	;
					tdata_save	[	30	]	<=	tdata_save	[	29	]	;
					tdata_save	[	31	]	<=	tdata_save	[	30	]	;
					tdata_save	[	32	]	<=	tdata_save	[	31	]	;
					tdata_save	[	33	]	<=	tdata_save	[	32	]	;
					tdata_save	[	34	]	<=	tdata_save	[	33	]	;
					tdata_save	[	35	]	<=	tdata_save	[	34	]	;
					tdata_save	[	36	]	<=	tdata_save	[	35	]	;
					tdata_save	[	37	]	<=	tdata_save	[	36	]	;
					tdata_save	[	38	]	<=	tdata_save	[	37	]	;
					tdata_save	[	39	]	<=	tdata_save	[	38	]	;
					tdata_save	[	40	]	<=	tdata_save	[	39	]	;
					tdata_save	[	41	]	<=	tdata_save	[	40	]	;
					tdata_save	[	42	]	<=	tdata_save	[	41	]	;
					tdata_save	[	43	]	<=	tdata_save	[	42	]	;
					tdata_save	[	44	]	<=	tdata_save	[	43	]	;
					tdata_save	[	45	]	<=	tdata_save	[	44	]	;
					tdata_save	[	46	]	<=	tdata_save	[	45	]	;
					tdata_save	[	47	]	<=	tdata_save	[	46	]	;
					tdata_save	[	48	]	<=	tdata_save	[	47	]	;
					tdata_save	[	49	]	<=	tdata_save	[	48	]	;
					tdata_save	[	50	]	<=	tdata_save	[	49	]	;
					tdata_save	[	51	]	<=	tdata_save	[	50	]	;
					tdata_save	[	52	]	<=	tdata_save	[	51	]	;
					tdata_save	[	53	]	<=	tdata_save	[	52	]	;
					tdata_save	[	54	]	<=	tdata_save	[	53	]	;
					tdata_save	[	55	]	<=	tdata_save	[	54	]	;
					tdata_save	[	56	]	<=	tdata_save	[	55	]	;
					tdata_save	[	57	]	<=	tdata_save	[	56	]	;
					tdata_save	[	58	]	<=	tdata_save	[	57	]	;
					tdata_save	[	59	]	<=	tdata_save	[	58	]	;
					tdata_save	[	60	]	<=	tdata_save	[	59	]	;
					tdata_save	[	61	]	<=	tdata_save	[	60	]	;
					tdata_save	[	62	]	<=	tdata_save	[	61	]	;
					tdata_save	[	63	]	<=	tdata_save	[	62	]	;
					tdata_save	[	64	]	<=	tdata_save	[	63	]	;
					tdata_save	[	65	]	<=	tdata_save	[	64	]	;
					tdata_save	[	66	]	<=	tdata_save	[	65	]	;
					tdata_save	[	67	]	<=	tdata_save	[	66	]	;
					tdata_save	[	68	]	<=	tdata_save	[	67	]	;
					tdata_save	[	69	]	<=	tdata_save	[	68	]	;
					tdata_save	[	70	]	<=	tdata_save	[	69	]	;
					tdata_save	[	71	]	<=	tdata_save	[	70	]	;
					tdata_save	[	72	]	<=	tdata_save	[	71	]	;
					tdata_save	[	73	]	<=	tdata_save	[	72	]	;
					tdata_save	[	74	]	<=	tdata_save	[	73	]	;
					tdata_save	[	75	]	<=	tdata_save	[	74	]	;
					tdata_save	[	76	]	<=	tdata_save	[	75	]	;
					tdata_save	[	77	]	<=	tdata_save	[	76	]	;
					tdata_save	[	78	]	<=	tdata_save	[	77	]	;
					tdata_save	[	79	]	<=	tdata_save	[	78	]	;
					tdata_save	[	80	]	<=	tdata_save	[	79	]	;
					tdata_save	[	81	]	<=	tdata_save	[	80	]	;
					tdata_save	[	82	]	<=	tdata_save	[	81	]	;
					tdata_save	[	83	]	<=	tdata_save	[	82	]	;
					tdata_save	[	84	]	<=	tdata_save	[	83	]	;
					tdata_save	[	85	]	<=	tdata_save	[	84	]	;
					tdata_save	[	86	]	<=	tdata_save	[	85	]	;
					tdata_save	[	87	]	<=	tdata_save	[	86	]	;
					tdata_save	[	88	]	<=	tdata_save	[	87	]	;
					tdata_save	[	89	]	<=	tdata_save	[	88	]	;
					tdata_save	[	90	]	<=	tdata_save	[	89	]	;
					tdata_save	[	91	]	<=	tdata_save	[	90	]	;
					tdata_save	[	92	]	<=	tdata_save	[	91	]	;
					tdata_save	[	93	]	<=	tdata_save	[	92	]	;
					tdata_save	[	94	]	<=	tdata_save	[	93	]	;
					tdata_save	[	95	]	<=	tdata_save	[	94	]	;
					tdata_save	[	96	]	<=	tdata_save	[	95	]	;
					tdata_save	[	97	]	<=	tdata_save	[	96	]	;
					tdata_save	[	98	]	<=	tdata_save	[	97	]	;
					tdata_save	[	99	]	<=	tdata_save	[	98	]	;
					tdata_save	[	100	]	<=	tdata_save	[	99	]	;
					tdata_save	[	101	]	<=	tdata_save	[	100	]	;
					tdata_save	[	102	]	<=	tdata_save	[	101	]	;
					tdata_save	[	103	]	<=	tdata_save	[	102	]	;
					tdata_save	[	104	]	<=	tdata_save	[	103	]	;
					tdata_save	[	105	]	<=	tdata_save	[	104	]	;
					tdata_save	[	106	]	<=	tdata_save	[	105	]	;
					tdata_save	[	107	]	<=	tdata_save	[	106	]	;
					tdata_save	[	108	]	<=	tdata_save	[	107	]	;
					tdata_save	[	109	]	<=	tdata_save	[	108	]	;
					tdata_save	[	110	]	<=	tdata_save	[	109	]	;
					tdata_save	[	111	]	<=	tdata_save	[	110	]	;
					tdata_save	[	112	]	<=	tdata_save	[	111	]	;
					tdata_save	[	113	]	<=	tdata_save	[	112	]	;
					tdata_save	[	114	]	<=	tdata_save	[	113	]	;
					tdata_save	[	115	]	<=	tdata_save	[	114	]	;
					tdata_save	[	116	]	<=	tdata_save	[	115	]	;
					tdata_save	[	117	]	<=	tdata_save	[	116	]	;
					tdata_save	[	118	]	<=	tdata_save	[	117	]	;
					tdata_save	[	119	]	<=	tdata_save	[	118	]	;
					tdata_save	[	120	]	<=	tdata_save	[	119	]	;
					tdata_save	[	121	]	<=	tdata_save	[	120	]	;
					tdata_save	[	122	]	<=	tdata_save	[	121	]	;
					tdata_save	[	123	]	<=	tdata_save	[	122	]	;
					tdata_save	[	124	]	<=	tdata_save	[	123	]	;
					tdata_save	[	125	]	<=	tdata_save	[	124	]	;
					tdata_save	[	126	]	<=	tdata_save	[	125	]	;
					tdata_save	[	127	]	<=	tdata_save	[	126	]	;
					tdata_save	[	128	]	<=	tdata_save	[	127	]	;
					tdata_save	[	129	]	<=	tdata_save	[	128	]	;
					tdata_save	[	130	]	<=	tdata_save	[	129	]	;
					tdata_save	[	131	]	<=	tdata_save	[	130	]	;
					tdata_save	[	132	]	<=	tdata_save	[	131	]	;
					tdata_save	[	133	]	<=	tdata_save	[	132	]	;
					tdata_save	[	134	]	<=	tdata_save	[	133	]	;
					tdata_save	[	135	]	<=	tdata_save	[	134	]	;
					tdata_save	[	136	]	<=	tdata_save	[	135	]	;
					tdata_save	[	137	]	<=	tdata_save	[	136	]	;
					tdata_save	[	138	]	<=	tdata_save	[	137	]	;
					tdata_save	[	139	]	<=	tdata_save	[	138	]	;
					tdata_save	[	140	]	<=	tdata_save	[	139	]	;
					tdata_save	[	141	]	<=	tdata_save	[	140	]	;
					tdata_save	[	142	]	<=	tdata_save	[	141	]	;
					tdata_save	[	143	]	<=	tdata_save	[	142	]	;
					tdata_save	[	144	]	<=	tdata_save	[	143	]	;
					tdata_save	[	145	]	<=	tdata_save	[	144	]	;
					tdata_save	[	146	]	<=	tdata_save	[	145	]	;
					tdata_save	[	147	]	<=	tdata_save	[	146	]	;
					tdata_save	[	148	]	<=	tdata_save	[	147	]	;
					tdata_save	[	149	]	<=	tdata_save	[	148	]	;
					tdata_save	[	150	]	<=	tdata_save	[	149	]	;
					tdata_save	[	151	]	<=	tdata_save	[	150	]	;
					tdata_save	[	152	]	<=	tdata_save	[	151	]	;
					tdata_save	[	153	]	<=	tdata_save	[	152	]	;
					tdata_save	[	154	]	<=	tdata_save	[	153	]	;
					tdata_save	[	155	]	<=	tdata_save	[	154	]	;
					tdata_save	[	156	]	<=	tdata_save	[	155	]	;
					tdata_save	[	157	]	<=	tdata_save	[	156	]	;
					tdata_save	[	158	]	<=	tdata_save	[	157	]	;
					tdata_save	[	159	]	<=	tdata_save	[	158	]	;
					tdata_save	[	160	]	<=	tdata_save	[	159	]	;
					tdata_save	[	161	]	<=	tdata_save	[	160	]	;
					tdata_save	[	162	]	<=	tdata_save	[	161	]	;
					tdata_save	[	163	]	<=	tdata_save	[	162	]	;
					tdata_save	[	164	]	<=	tdata_save	[	163	]	;
					tdata_save	[	165	]	<=	tdata_save	[	164	]	;
					tdata_save	[	166	]	<=	tdata_save	[	165	]	;
					tdata_save	[	167	]	<=	tdata_save	[	166	]	;
					tdata_save	[	168	]	<=	tdata_save	[	167	]	;
					tdata_save	[	169	]	<=	tdata_save	[	168	]	;
					tdata_save	[	170	]	<=	tdata_save	[	169	]	;
					tdata_save	[	171	]	<=	tdata_save	[	170	]	;
					tdata_save	[	172	]	<=	tdata_save	[	171	]	;
					tdata_save	[	173	]	<=	tdata_save	[	172	]	;
					tdata_save	[	174	]	<=	tdata_save	[	173	]	;
					tdata_save	[	175	]	<=	tdata_save	[	174	]	;
					tdata_save	[	176	]	<=	tdata_save	[	175	]	;
					tdata_save	[	177	]	<=	tdata_save	[	176	]	;
					tdata_save	[	178	]	<=	tdata_save	[	177	]	;
					tdata_save	[	179	]	<=	tdata_save	[	178	]	;
					tdata_save	[	180	]	<=	tdata_save	[	179	]	;
					tdata_save	[	181	]	<=	tdata_save	[	180	]	;
					tdata_save	[	182	]	<=	tdata_save	[	181	]	;
					tdata_save	[	183	]	<=	tdata_save	[	182	]	;
					tdata_save	[	184	]	<=	tdata_save	[	183	]	;
					tdata_save	[	185	]	<=	tdata_save	[	184	]	;
					tdata_save	[	186	]	<=	tdata_save	[	185	]	;
					tdata_save	[	187	]	<=	tdata_save	[	186	]	;
					tdata_save	[	188	]	<=	tdata_save	[	187	]	;
					tdata_save	[	189	]	<=	tdata_save	[	188	]	;
					tdata_save	[	190	]	<=	tdata_save	[	189	]	;
					tdata_save	[	191	]	<=	tdata_save	[	190	]	;
					tdata_save	[	192	]	<=	tdata_save	[	191	]	;
					tdata_save	[	193	]	<=	tdata_save	[	192	]	;
					tdata_save	[	194	]	<=	tdata_save	[	193	]	;
					tdata_save	[	195	]	<=	tdata_save	[	194	]	;
					tdata_save	[	196	]	<=	tdata_save	[	195	]	;
					tdata_save	[	197	]	<=	tdata_save	[	196	]	;
					tdata_save	[	198	]	<=	tdata_save	[	197	]	;
					tdata_save	[	199	]	<=	tdata_save	[	198	]	;
					tdata_save	[	200	]	<=	tdata_save	[	199	]	;
					tdata_save	[	201	]	<=	tdata_save	[	200	]	;
					tdata_save	[	202	]	<=	tdata_save	[	201	]	;
					tdata_save	[	203	]	<=	tdata_save	[	202	]	;
					tdata_save	[	204	]	<=	tdata_save	[	203	]	;
					tdata_save	[	205	]	<=	tdata_save	[	204	]	;
					tdata_save	[	206	]	<=	tdata_save	[	205	]	;
					tdata_save	[	207	]	<=	tdata_save	[	206	]	;
					tdata_save	[	208	]	<=	tdata_save	[	207	]	;
					tdata_save	[	209	]	<=	tdata_save	[	208	]	;
					tdata_save	[	210	]	<=	tdata_save	[	209	]	;
					tdata_save	[	211	]	<=	tdata_save	[	210	]	;
					tdata_save	[	212	]	<=	tdata_save	[	211	]	;
					tdata_save	[	213	]	<=	tdata_save	[	212	]	;
					tdata_save	[	214	]	<=	tdata_save	[	213	]	;
					tdata_save	[	215	]	<=	tdata_save	[	214	]	;
					tdata_save	[	216	]	<=	tdata_save	[	215	]	;
					tdata_save	[	217	]	<=	tdata_save	[	216	]	;
					tdata_save	[	218	]	<=	tdata_save	[	217	]	;
					tdata_save	[	219	]	<=	tdata_save	[	218	]	;
					tdata_save	[	220	]	<=	tdata_save	[	219	]	;
					tdata_save	[	221	]	<=	tdata_save	[	220	]	;
					tdata_save	[	222	]	<=	tdata_save	[	221	]	;
					tdata_save	[	223	]	<=	tdata_save	[	222	]	;
					tdata_save	[	224	]	<=	tdata_save	[	223	]	;
					tdata_save	[	225	]	<=	tdata_save	[	224	]	;
					tdata_save	[	226	]	<=	tdata_save	[	225	]	;
					tdata_save	[	227	]	<=	tdata_save	[	226	]	;
					tdata_save	[	228	]	<=	tdata_save	[	227	]	;
					tdata_save	[	229	]	<=	tdata_save	[	228	]	;
					tdata_save	[	230	]	<=	tdata_save	[	229	]	;
					tdata_save	[	231	]	<=	tdata_save	[	230	]	;
					tdata_save	[	232	]	<=	tdata_save	[	231	]	;
					tdata_save	[	233	]	<=	tdata_save	[	232	]	;
					tdata_save	[	234	]	<=	tdata_save	[	233	]	;
					tdata_save	[	235	]	<=	tdata_save	[	234	]	;
					tdata_save	[	236	]	<=	tdata_save	[	235	]	;
					tdata_save	[	237	]	<=	tdata_save	[	236	]	;
					tdata_save	[	238	]	<=	tdata_save	[	237	]	;
					tdata_save	[	239	]	<=	tdata_save	[	238	]	;
					tdata_save	[	240	]	<=	tdata_save	[	239	]	;
					tdata_save	[	241	]	<=	tdata_save	[	240	]	;
					tdata_save	[	242	]	<=	tdata_save	[	241	]	;
					tdata_save	[	243	]	<=	tdata_save	[	242	]	;
					tdata_save	[	244	]	<=	tdata_save	[	243	]	;
					tdata_save	[	245	]	<=	tdata_save	[	244	]	;
					tdata_save	[	246	]	<=	tdata_save	[	245	]	;
					tdata_save	[	247	]	<=	tdata_save	[	246	]	;
					tdata_save	[	248	]	<=	tdata_save	[	247	]	;
					tdata_save	[	249	]	<=	tdata_save	[	248	]	;
					tdata_save	[	250	]	<=	tdata_save	[	249	]	;
					tdata_save	[	251	]	<=	tdata_save	[	250	]	;
					tdata_save	[	252	]	<=	tdata_save	[	251	]	;
					tdata_save	[	253	]	<=	tdata_save	[	252	]	;
					tdata_save	[	254	]	<=	tdata_save	[	253	]	;
					tdata_save	[	255	]	<=	tdata_save	[	254	]	;
					tuser_save	[	0	]	<=	tuser;						
				tuser_save	[	1	]	<=	tuser_save	[	0	]	;
				tuser_save	[	2	]	<=	tuser_save	[	1	]	;
				tuser_save	[	3	]	<=	tuser_save	[	2	]	;
				tuser_save	[	4	]	<=	tuser_save	[	3	]	;
				tuser_save	[	5	]	<=	tuser_save	[	4	]	;
				tuser_save	[	6	]	<=	tuser_save	[	5	]	;
				tuser_save	[	7	]	<=	tuser_save	[	6	]	;
				tuser_save	[	8	]	<=	tuser_save	[	7	]	;
				tuser_save	[	9	]	<=	tuser_save	[	8	]	;
				tuser_save	[	10	]	<=	tuser_save	[	9	]	;
				tuser_save	[	11	]	<=	tuser_save	[	10	]	;
				tuser_save	[	12	]	<=	tuser_save	[	11	]	;
				tuser_save	[	13	]	<=	tuser_save	[	12	]	;
				tuser_save	[	14	]	<=	tuser_save	[	13	]	;
				tuser_save	[	15	]	<=	tuser_save	[	14	]	;
				tuser_save	[	16	]	<=	tuser_save	[	15	]	;
				tuser_save	[	17	]	<=	tuser_save	[	16	]	;
				tuser_save	[	18	]	<=	tuser_save	[	17	]	;
				tuser_save	[	19	]	<=	tuser_save	[	18	]	;
				tuser_save	[	20	]	<=	tuser_save	[	19	]	;
				tuser_save	[	21	]	<=	tuser_save	[	20	]	;
				tuser_save	[	22	]	<=	tuser_save	[	21	]	;
				tuser_save	[	23	]	<=	tuser_save	[	22	]	;
				tuser_save	[	24	]	<=	tuser_save	[	23	]	;
				tuser_save	[	25	]	<=	tuser_save	[	24	]	;
				tuser_save	[	26	]	<=	tuser_save	[	25	]	;
				tuser_save	[	27	]	<=	tuser_save	[	26	]	;
				tuser_save	[	28	]	<=	tuser_save	[	27	]	;
				tuser_save	[	29	]	<=	tuser_save	[	28	]	;
				tuser_save	[	30	]	<=	tuser_save	[	29	]	;
				tuser_save	[	31	]	<=	tuser_save	[	30	]	;
				tuser_save	[	32	]	<=	tuser_save	[	31	]	;
				tuser_save	[	33	]	<=	tuser_save	[	32	]	;
				tuser_save	[	34	]	<=	tuser_save	[	33	]	;
				tuser_save	[	35	]	<=	tuser_save	[	34	]	;
				tuser_save	[	36	]	<=	tuser_save	[	35	]	;
				tuser_save	[	37	]	<=	tuser_save	[	36	]	;
				tuser_save	[	38	]	<=	tuser_save	[	37	]	;
				tuser_save	[	39	]	<=	tuser_save	[	38	]	;
				tuser_save	[	40	]	<=	tuser_save	[	39	]	;
				tuser_save	[	41	]	<=	tuser_save	[	40	]	;
				tuser_save	[	42	]	<=	tuser_save	[	41	]	;
				tuser_save	[	43	]	<=	tuser_save	[	42	]	;
				tuser_save	[	44	]	<=	tuser_save	[	43	]	;
				tuser_save	[	45	]	<=	tuser_save	[	44	]	;
				tuser_save	[	46	]	<=	tuser_save	[	45	]	;
				tuser_save	[	47	]	<=	tuser_save	[	46	]	;
				tuser_save	[	48	]	<=	tuser_save	[	47	]	;
				tuser_save	[	49	]	<=	tuser_save	[	48	]	;
				tuser_save	[	50	]	<=	tuser_save	[	49	]	;
				tuser_save	[	51	]	<=	tuser_save	[	50	]	;
				tuser_save	[	52	]	<=	tuser_save	[	51	]	;
				tuser_save	[	53	]	<=	tuser_save	[	52	]	;
				tuser_save	[	54	]	<=	tuser_save	[	53	]	;
				tuser_save	[	55	]	<=	tuser_save	[	54	]	;
				tuser_save	[	56	]	<=	tuser_save	[	55	]	;
				tuser_save	[	57	]	<=	tuser_save	[	56	]	;
				tuser_save	[	58	]	<=	tuser_save	[	57	]	;
				tuser_save	[	59	]	<=	tuser_save	[	58	]	;
				tuser_save	[	60	]	<=	tuser_save	[	59	]	;
				tuser_save	[	61	]	<=	tuser_save	[	60	]	;
				tuser_save	[	62	]	<=	tuser_save	[	61	]	;
				tuser_save	[	63	]	<=	tuser_save	[	62	]	;
				tuser_save	[	64	]	<=	tuser_save	[	63	]	;
				tuser_save	[	65	]	<=	tuser_save	[	64	]	;
				tuser_save	[	66	]	<=	tuser_save	[	65	]	;
				tuser_save	[	67	]	<=	tuser_save	[	66	]	;
				tuser_save	[	68	]	<=	tuser_save	[	67	]	;
				tuser_save	[	69	]	<=	tuser_save	[	68	]	;
				tuser_save	[	70	]	<=	tuser_save	[	69	]	;
				tuser_save	[	71	]	<=	tuser_save	[	70	]	;
				tuser_save	[	72	]	<=	tuser_save	[	71	]	;
				tuser_save	[	73	]	<=	tuser_save	[	72	]	;
				tuser_save	[	74	]	<=	tuser_save	[	73	]	;
				tuser_save	[	75	]	<=	tuser_save	[	74	]	;
				tuser_save	[	76	]	<=	tuser_save	[	75	]	;
				tuser_save	[	77	]	<=	tuser_save	[	76	]	;
				tuser_save	[	78	]	<=	tuser_save	[	77	]	;
				tuser_save	[	79	]	<=	tuser_save	[	78	]	;
				tuser_save	[	80	]	<=	tuser_save	[	79	]	;
				tuser_save	[	81	]	<=	tuser_save	[	80	]	;
				tuser_save	[	82	]	<=	tuser_save	[	81	]	;
				tuser_save	[	83	]	<=	tuser_save	[	82	]	;
				tuser_save	[	84	]	<=	tuser_save	[	83	]	;
				tuser_save	[	85	]	<=	tuser_save	[	84	]	;
				tuser_save	[	86	]	<=	tuser_save	[	85	]	;
				tuser_save	[	87	]	<=	tuser_save	[	86	]	;
				tuser_save	[	88	]	<=	tuser_save	[	87	]	;
				tuser_save	[	89	]	<=	tuser_save	[	88	]	;
				tuser_save	[	90	]	<=	tuser_save	[	89	]	;
				tuser_save	[	91	]	<=	tuser_save	[	90	]	;
				tuser_save	[	92	]	<=	tuser_save	[	91	]	;
				tuser_save	[	93	]	<=	tuser_save	[	92	]	;
				tuser_save	[	94	]	<=	tuser_save	[	93	]	;
				tuser_save	[	95	]	<=	tuser_save	[	94	]	;
				tuser_save	[	96	]	<=	tuser_save	[	95	]	;
				tuser_save	[	97	]	<=	tuser_save	[	96	]	;
				tuser_save	[	98	]	<=	tuser_save	[	97	]	;
				tuser_save	[	99	]	<=	tuser_save	[	98	]	;
				tuser_save	[	100	]	<=	tuser_save	[	99	]	;
				tuser_save	[	101	]	<=	tuser_save	[	100	]	;
				tuser_save	[	102	]	<=	tuser_save	[	101	]	;
				tuser_save	[	103	]	<=	tuser_save	[	102	]	;
				tuser_save	[	104	]	<=	tuser_save	[	103	]	;
				tuser_save	[	105	]	<=	tuser_save	[	104	]	;
				tuser_save	[	106	]	<=	tuser_save	[	105	]	;
				tuser_save	[	107	]	<=	tuser_save	[	106	]	;
				tuser_save	[	108	]	<=	tuser_save	[	107	]	;
				tuser_save	[	109	]	<=	tuser_save	[	108	]	;
				tuser_save	[	110	]	<=	tuser_save	[	109	]	;
				tuser_save	[	111	]	<=	tuser_save	[	110	]	;
				tuser_save	[	112	]	<=	tuser_save	[	111	]	;
				tuser_save	[	113	]	<=	tuser_save	[	112	]	;
				tuser_save	[	114	]	<=	tuser_save	[	113	]	;
				tuser_save	[	115	]	<=	tuser_save	[	114	]	;
				tuser_save	[	116	]	<=	tuser_save	[	115	]	;
				tuser_save	[	117	]	<=	tuser_save	[	116	]	;
				tuser_save	[	118	]	<=	tuser_save	[	117	]	;
				tuser_save	[	119	]	<=	tuser_save	[	118	]	;
				tuser_save	[	120	]	<=	tuser_save	[	119	]	;
				tuser_save	[	121	]	<=	tuser_save	[	120	]	;
				tuser_save	[	122	]	<=	tuser_save	[	121	]	;
				tuser_save	[	123	]	<=	tuser_save	[	122	]	;
				tuser_save	[	124	]	<=	tuser_save	[	123	]	;
				tuser_save	[	125	]	<=	tuser_save	[	124	]	;
				tuser_save	[	126	]	<=	tuser_save	[	125	]	;
				tuser_save	[	127	]	<=	tuser_save	[	126	]	;
				tuser_save	[	128	]	<=	tuser_save	[	127	]	;
				tuser_save	[	129	]	<=	tuser_save	[	128	]	;
				tuser_save	[	130	]	<=	tuser_save	[	129	]	;
				tuser_save	[	131	]	<=	tuser_save	[	130	]	;
				tuser_save	[	132	]	<=	tuser_save	[	131	]	;
				tuser_save	[	133	]	<=	tuser_save	[	132	]	;
				tuser_save	[	134	]	<=	tuser_save	[	133	]	;
				tuser_save	[	135	]	<=	tuser_save	[	134	]	;
				tuser_save	[	136	]	<=	tuser_save	[	135	]	;
				tuser_save	[	137	]	<=	tuser_save	[	136	]	;
				tuser_save	[	138	]	<=	tuser_save	[	137	]	;
				tuser_save	[	139	]	<=	tuser_save	[	138	]	;
				tuser_save	[	140	]	<=	tuser_save	[	139	]	;
				tuser_save	[	141	]	<=	tuser_save	[	140	]	;
				tuser_save	[	142	]	<=	tuser_save	[	141	]	;
				tuser_save	[	143	]	<=	tuser_save	[	142	]	;
				tuser_save	[	144	]	<=	tuser_save	[	143	]	;
				tuser_save	[	145	]	<=	tuser_save	[	144	]	;
				tuser_save	[	146	]	<=	tuser_save	[	145	]	;
				tuser_save	[	147	]	<=	tuser_save	[	146	]	;
				tuser_save	[	148	]	<=	tuser_save	[	147	]	;
				tuser_save	[	149	]	<=	tuser_save	[	148	]	;
				tuser_save	[	150	]	<=	tuser_save	[	149	]	;
				tuser_save	[	151	]	<=	tuser_save	[	150	]	;
				tuser_save	[	152	]	<=	tuser_save	[	151	]	;
				tuser_save	[	153	]	<=	tuser_save	[	152	]	;
				tuser_save	[	154	]	<=	tuser_save	[	153	]	;
				tuser_save	[	155	]	<=	tuser_save	[	154	]	;
				tuser_save	[	156	]	<=	tuser_save	[	155	]	;
				tuser_save	[	157	]	<=	tuser_save	[	156	]	;
				tuser_save	[	158	]	<=	tuser_save	[	157	]	;
				tuser_save	[	159	]	<=	tuser_save	[	158	]	;
				tuser_save	[	160	]	<=	tuser_save	[	159	]	;
				tuser_save	[	161	]	<=	tuser_save	[	160	]	;
				tuser_save	[	162	]	<=	tuser_save	[	161	]	;
				tuser_save	[	163	]	<=	tuser_save	[	162	]	;
				tuser_save	[	164	]	<=	tuser_save	[	163	]	;
				tuser_save	[	165	]	<=	tuser_save	[	164	]	;
				tuser_save	[	166	]	<=	tuser_save	[	165	]	;
				tuser_save	[	167	]	<=	tuser_save	[	166	]	;
				tuser_save	[	168	]	<=	tuser_save	[	167	]	;
				tuser_save	[	169	]	<=	tuser_save	[	168	]	;
				tuser_save	[	170	]	<=	tuser_save	[	169	]	;
				tuser_save	[	171	]	<=	tuser_save	[	170	]	;
				tuser_save	[	172	]	<=	tuser_save	[	171	]	;
				tuser_save	[	173	]	<=	tuser_save	[	172	]	;
				tuser_save	[	174	]	<=	tuser_save	[	173	]	;
				tuser_save	[	175	]	<=	tuser_save	[	174	]	;
				tuser_save	[	176	]	<=	tuser_save	[	175	]	;
				tuser_save	[	177	]	<=	tuser_save	[	176	]	;
				tuser_save	[	178	]	<=	tuser_save	[	177	]	;
				tuser_save	[	179	]	<=	tuser_save	[	178	]	;
				tuser_save	[	180	]	<=	tuser_save	[	179	]	;
				tuser_save	[	181	]	<=	tuser_save	[	180	]	;
				tuser_save	[	182	]	<=	tuser_save	[	181	]	;
				tuser_save	[	183	]	<=	tuser_save	[	182	]	;
				tuser_save	[	184	]	<=	tuser_save	[	183	]	;
				tuser_save	[	185	]	<=	tuser_save	[	184	]	;
				tuser_save	[	186	]	<=	tuser_save	[	185	]	;
				tuser_save	[	187	]	<=	tuser_save	[	186	]	;
				tuser_save	[	188	]	<=	tuser_save	[	187	]	;
				tuser_save	[	189	]	<=	tuser_save	[	188	]	;
				tuser_save	[	190	]	<=	tuser_save	[	189	]	;
				tuser_save	[	191	]	<=	tuser_save	[	190	]	;
				tuser_save	[	192	]	<=	tuser_save	[	191	]	;
				tuser_save	[	193	]	<=	tuser_save	[	192	]	;
				tuser_save	[	194	]	<=	tuser_save	[	193	]	;
				tuser_save	[	195	]	<=	tuser_save	[	194	]	;
				tuser_save	[	196	]	<=	tuser_save	[	195	]	;
				tuser_save	[	197	]	<=	tuser_save	[	196	]	;
				tuser_save	[	198	]	<=	tuser_save	[	197	]	;
				tuser_save	[	199	]	<=	tuser_save	[	198	]	;
				tuser_save	[	200	]	<=	tuser_save	[	199	]	;
				tuser_save	[	201	]	<=	tuser_save	[	200	]	;
				tuser_save	[	202	]	<=	tuser_save	[	201	]	;
				tuser_save	[	203	]	<=	tuser_save	[	202	]	;
				tuser_save	[	204	]	<=	tuser_save	[	203	]	;
				tuser_save	[	205	]	<=	tuser_save	[	204	]	;
				tuser_save	[	206	]	<=	tuser_save	[	205	]	;
				tuser_save	[	207	]	<=	tuser_save	[	206	]	;
				tuser_save	[	208	]	<=	tuser_save	[	207	]	;
				tuser_save	[	209	]	<=	tuser_save	[	208	]	;
				tuser_save	[	210	]	<=	tuser_save	[	209	]	;
				tuser_save	[	211	]	<=	tuser_save	[	210	]	;
				tuser_save	[	212	]	<=	tuser_save	[	211	]	;
				tuser_save	[	213	]	<=	tuser_save	[	212	]	;
				tuser_save	[	214	]	<=	tuser_save	[	213	]	;
				tuser_save	[	215	]	<=	tuser_save	[	214	]	;
				tuser_save	[	216	]	<=	tuser_save	[	215	]	;
				tuser_save	[	217	]	<=	tuser_save	[	216	]	;
				tuser_save	[	218	]	<=	tuser_save	[	217	]	;
				tuser_save	[	219	]	<=	tuser_save	[	218	]	;
				tuser_save	[	220	]	<=	tuser_save	[	219	]	;
				tuser_save	[	221	]	<=	tuser_save	[	220	]	;
				tuser_save	[	222	]	<=	tuser_save	[	221	]	;
				tuser_save	[	223	]	<=	tuser_save	[	222	]	;
				tuser_save	[	224	]	<=	tuser_save	[	223	]	;
				tuser_save	[	225	]	<=	tuser_save	[	224	]	;
				tuser_save	[	226	]	<=	tuser_save	[	225	]	;
				tuser_save	[	227	]	<=	tuser_save	[	226	]	;
				tuser_save	[	228	]	<=	tuser_save	[	227	]	;
				tuser_save	[	229	]	<=	tuser_save	[	228	]	;
				tuser_save	[	230	]	<=	tuser_save	[	229	]	;
				tuser_save	[	231	]	<=	tuser_save	[	230	]	;
				tuser_save	[	232	]	<=	tuser_save	[	231	]	;
				tuser_save	[	233	]	<=	tuser_save	[	232	]	;
				tuser_save	[	234	]	<=	tuser_save	[	233	]	;
				tuser_save	[	235	]	<=	tuser_save	[	234	]	;
				tuser_save	[	236	]	<=	tuser_save	[	235	]	;
				tuser_save	[	237	]	<=	tuser_save	[	236	]	;
				tuser_save	[	238	]	<=	tuser_save	[	237	]	;
				tuser_save	[	239	]	<=	tuser_save	[	238	]	;
				tuser_save	[	240	]	<=	tuser_save	[	239	]	;
				tuser_save	[	241	]	<=	tuser_save	[	240	]	;
				tuser_save	[	242	]	<=	tuser_save	[	241	]	;
				tuser_save	[	243	]	<=	tuser_save	[	242	]	;
				tuser_save	[	244	]	<=	tuser_save	[	243	]	;
				tuser_save	[	245	]	<=	tuser_save	[	244	]	;
				tuser_save	[	246	]	<=	tuser_save	[	245	]	;
				tuser_save	[	247	]	<=	tuser_save	[	246	]	;
				tuser_save	[	248	]	<=	tuser_save	[	247	]	;
				tuser_save	[	249	]	<=	tuser_save	[	248	]	;
				tuser_save	[	250	]	<=	tuser_save	[	249	]	;
				tuser_save	[	251	]	<=	tuser_save	[	250	]	;
				tuser_save	[	252	]	<=	tuser_save	[	251	]	;
				tuser_save	[	253	]	<=	tuser_save	[	252	]	;
				tuser_save	[	254	]	<=	tuser_save	[	253	]	;
				tuser_save	[	255	]	<=	tuser_save	[	254	]	;
					if(count_packet == 2'd2)
					begin
						count_packet <= 2'd0;
					end
					else
					begin
						count_packet	<= count_packet + 1'b1;
					end
					sum_tdata		<=	201'd0;
					sum_tuser		<=	128'd0;
					sum_tdata_valid		<=	1'b0;
					sum_tuser_valid		<=	1'b0;
				end
				else
				begin
					tdata_save	[	0	]	<=	tdata_save	[	0	]	;//stay_no_change
					tdata_save	[	1	]	<=	tdata_save	[	1	]	;
					tdata_save	[	2	]	<=	tdata_save	[	2	]	;
					tdata_save	[	3	]	<=	tdata_save	[	3	]	;
					tdata_save	[	4	]	<=	tdata_save	[	4	]	;
					tdata_save	[	5	]	<=	tdata_save	[	5	]	;
					tdata_save	[	6	]	<=	tdata_save	[	6	]	;
					tdata_save	[	7	]	<=	tdata_save	[	7	]	;
					tdata_save	[	8	]	<=	tdata_save	[	8	]	;
					tdata_save	[	9	]	<=	tdata_save	[	9	]	;
					tdata_save	[	10	]	<=	tdata_save	[	10	]	;
					tdata_save	[	11	]	<=	tdata_save	[	11	]	;
					tdata_save	[	12	]	<=	tdata_save	[	12	]	;
					tdata_save	[	13	]	<=	tdata_save	[	13	]	;
					tdata_save	[	14	]	<=	tdata_save	[	14	]	;
					tdata_save	[	15	]	<=	tdata_save	[	15	]	;
					tdata_save	[	16	]	<=	tdata_save	[	16	]	;
					tdata_save	[	17	]	<=	tdata_save	[	17	]	;
					tdata_save	[	18	]	<=	tdata_save	[	18	]	;
					tdata_save	[	19	]	<=	tdata_save	[	19	]	;
					tdata_save	[	20	]	<=	tdata_save	[	20	]	;
					tdata_save	[	21	]	<=	tdata_save	[	21	]	;
					tdata_save	[	22	]	<=	tdata_save	[	22	]	;
					tdata_save	[	23	]	<=	tdata_save	[	23	]	;
					tdata_save	[	24	]	<=	tdata_save	[	24	]	;
					tdata_save	[	25	]	<=	tdata_save	[	25	]	;
					tdata_save	[	26	]	<=	tdata_save	[	26	]	;
					tdata_save	[	27	]	<=	tdata_save	[	27	]	;
					tdata_save	[	28	]	<=	tdata_save	[	28	]	;
					tdata_save	[	29	]	<=	tdata_save	[	29	]	;
					tdata_save	[	30	]	<=	tdata_save	[	30	]	;
					tdata_save	[	31	]	<=	tdata_save	[	31	]	;
					tdata_save	[	32	]	<=	tdata_save	[	32	]	;
					tdata_save	[	33	]	<=	tdata_save	[	33	]	;
					tdata_save	[	34	]	<=	tdata_save	[	34	]	;
					tdata_save	[	35	]	<=	tdata_save	[	35	]	;
					tdata_save	[	36	]	<=	tdata_save	[	36	]	;
					tdata_save	[	37	]	<=	tdata_save	[	37	]	;
					tdata_save	[	38	]	<=	tdata_save	[	38	]	;
					tdata_save	[	39	]	<=	tdata_save	[	39	]	;
					tdata_save	[	40	]	<=	tdata_save	[	40	]	;
					tdata_save	[	41	]	<=	tdata_save	[	41	]	;
					tdata_save	[	42	]	<=	tdata_save	[	42	]	;
					tdata_save	[	43	]	<=	tdata_save	[	43	]	;
					tdata_save	[	44	]	<=	tdata_save	[	44	]	;
					tdata_save	[	45	]	<=	tdata_save	[	45	]	;
					tdata_save	[	46	]	<=	tdata_save	[	46	]	;
					tdata_save	[	47	]	<=	tdata_save	[	47	]	;
					tdata_save	[	48	]	<=	tdata_save	[	48	]	;
					tdata_save	[	49	]	<=	tdata_save	[	49	]	;
					tdata_save	[	50	]	<=	tdata_save	[	50	]	;
					tdata_save	[	51	]	<=	tdata_save	[	51	]	;
					tdata_save	[	52	]	<=	tdata_save	[	52	]	;
					tdata_save	[	53	]	<=	tdata_save	[	53	]	;
					tdata_save	[	54	]	<=	tdata_save	[	54	]	;
					tdata_save	[	55	]	<=	tdata_save	[	55	]	;
					tdata_save	[	56	]	<=	tdata_save	[	56	]	;
					tdata_save	[	57	]	<=	tdata_save	[	57	]	;
					tdata_save	[	58	]	<=	tdata_save	[	58	]	;
					tdata_save	[	59	]	<=	tdata_save	[	59	]	;
					tdata_save	[	60	]	<=	tdata_save	[	60	]	;
					tdata_save	[	61	]	<=	tdata_save	[	61	]	;
					tdata_save	[	62	]	<=	tdata_save	[	62	]	;
					tdata_save	[	63	]	<=	tdata_save	[	63	]	;
					tdata_save	[	64	]	<=	tdata_save	[	64	]	;
					tdata_save	[	65	]	<=	tdata_save	[	65	]	;
					tdata_save	[	66	]	<=	tdata_save	[	66	]	;
					tdata_save	[	67	]	<=	tdata_save	[	67	]	;
					tdata_save	[	68	]	<=	tdata_save	[	68	]	;
					tdata_save	[	69	]	<=	tdata_save	[	69	]	;
					tdata_save	[	70	]	<=	tdata_save	[	70	]	;
					tdata_save	[	71	]	<=	tdata_save	[	71	]	;
					tdata_save	[	72	]	<=	tdata_save	[	72	]	;
					tdata_save	[	73	]	<=	tdata_save	[	73	]	;
					tdata_save	[	74	]	<=	tdata_save	[	74	]	;
					tdata_save	[	75	]	<=	tdata_save	[	75	]	;
					tdata_save	[	76	]	<=	tdata_save	[	76	]	;
					tdata_save	[	77	]	<=	tdata_save	[	77	]	;
					tdata_save	[	78	]	<=	tdata_save	[	78	]	;
					tdata_save	[	79	]	<=	tdata_save	[	79	]	;
					tdata_save	[	80	]	<=	tdata_save	[	80	]	;
					tdata_save	[	81	]	<=	tdata_save	[	81	]	;
					tdata_save	[	82	]	<=	tdata_save	[	82	]	;
					tdata_save	[	83	]	<=	tdata_save	[	83	]	;
					tdata_save	[	84	]	<=	tdata_save	[	84	]	;
					tdata_save	[	85	]	<=	tdata_save	[	85	]	;
					tdata_save	[	86	]	<=	tdata_save	[	86	]	;
					tdata_save	[	87	]	<=	tdata_save	[	87	]	;
					tdata_save	[	88	]	<=	tdata_save	[	88	]	;
					tdata_save	[	89	]	<=	tdata_save	[	89	]	;
					tdata_save	[	90	]	<=	tdata_save	[	90	]	;
					tdata_save	[	91	]	<=	tdata_save	[	91	]	;
					tdata_save	[	92	]	<=	tdata_save	[	92	]	;
					tdata_save	[	93	]	<=	tdata_save	[	93	]	;
					tdata_save	[	94	]	<=	tdata_save	[	94	]	;
					tdata_save	[	95	]	<=	tdata_save	[	95	]	;
					tdata_save	[	96	]	<=	tdata_save	[	96	]	;
					tdata_save	[	97	]	<=	tdata_save	[	97	]	;
					tdata_save	[	98	]	<=	tdata_save	[	98	]	;
					tdata_save	[	99	]	<=	tdata_save	[	99	]	;
					tdata_save	[	100	]	<=	tdata_save	[	100	]	;
					tdata_save	[	101	]	<=	tdata_save	[	101	]	;
					tdata_save	[	102	]	<=	tdata_save	[	102	]	;
					tdata_save	[	103	]	<=	tdata_save	[	103	]	;
					tdata_save	[	104	]	<=	tdata_save	[	104	]	;
					tdata_save	[	105	]	<=	tdata_save	[	105	]	;
					tdata_save	[	106	]	<=	tdata_save	[	106	]	;
					tdata_save	[	107	]	<=	tdata_save	[	107	]	;
					tdata_save	[	108	]	<=	tdata_save	[	108	]	;
					tdata_save	[	109	]	<=	tdata_save	[	109	]	;
					tdata_save	[	110	]	<=	tdata_save	[	110	]	;
					tdata_save	[	111	]	<=	tdata_save	[	111	]	;
					tdata_save	[	112	]	<=	tdata_save	[	112	]	;
					tdata_save	[	113	]	<=	tdata_save	[	113	]	;
					tdata_save	[	114	]	<=	tdata_save	[	114	]	;
					tdata_save	[	115	]	<=	tdata_save	[	115	]	;
					tdata_save	[	116	]	<=	tdata_save	[	116	]	;
					tdata_save	[	117	]	<=	tdata_save	[	117	]	;
					tdata_save	[	118	]	<=	tdata_save	[	118	]	;
					tdata_save	[	119	]	<=	tdata_save	[	119	]	;
					tdata_save	[	120	]	<=	tdata_save	[	120	]	;
					tdata_save	[	121	]	<=	tdata_save	[	121	]	;
					tdata_save	[	122	]	<=	tdata_save	[	122	]	;
					tdata_save	[	123	]	<=	tdata_save	[	123	]	;
					tdata_save	[	124	]	<=	tdata_save	[	124	]	;
					tdata_save	[	125	]	<=	tdata_save	[	125	]	;
					tdata_save	[	126	]	<=	tdata_save	[	126	]	;
					tdata_save	[	127	]	<=	tdata_save	[	127	]	;
					tdata_save	[	128	]	<=	tdata_save	[	128	]	;
					tdata_save	[	129	]	<=	tdata_save	[	129	]	;
					tdata_save	[	130	]	<=	tdata_save	[	130	]	;
					tdata_save	[	131	]	<=	tdata_save	[	131	]	;
					tdata_save	[	132	]	<=	tdata_save	[	132	]	;
					tdata_save	[	133	]	<=	tdata_save	[	133	]	;
					tdata_save	[	134	]	<=	tdata_save	[	134	]	;
					tdata_save	[	135	]	<=	tdata_save	[	135	]	;
					tdata_save	[	136	]	<=	tdata_save	[	136	]	;
					tdata_save	[	137	]	<=	tdata_save	[	137	]	;
					tdata_save	[	138	]	<=	tdata_save	[	138	]	;
					tdata_save	[	139	]	<=	tdata_save	[	139	]	;
					tdata_save	[	140	]	<=	tdata_save	[	140	]	;
					tdata_save	[	141	]	<=	tdata_save	[	141	]	;
					tdata_save	[	142	]	<=	tdata_save	[	142	]	;
					tdata_save	[	143	]	<=	tdata_save	[	143	]	;
					tdata_save	[	144	]	<=	tdata_save	[	144	]	;
					tdata_save	[	145	]	<=	tdata_save	[	145	]	;
					tdata_save	[	146	]	<=	tdata_save	[	146	]	;
					tdata_save	[	147	]	<=	tdata_save	[	147	]	;
					tdata_save	[	148	]	<=	tdata_save	[	148	]	;
					tdata_save	[	149	]	<=	tdata_save	[	149	]	;
					tdata_save	[	150	]	<=	tdata_save	[	150	]	;
					tdata_save	[	151	]	<=	tdata_save	[	151	]	;
					tdata_save	[	152	]	<=	tdata_save	[	152	]	;
					tdata_save	[	153	]	<=	tdata_save	[	153	]	;
					tdata_save	[	154	]	<=	tdata_save	[	154	]	;
					tdata_save	[	155	]	<=	tdata_save	[	155	]	;
					tdata_save	[	156	]	<=	tdata_save	[	156	]	;
					tdata_save	[	157	]	<=	tdata_save	[	157	]	;
					tdata_save	[	158	]	<=	tdata_save	[	158	]	;
					tdata_save	[	159	]	<=	tdata_save	[	159	]	;
					tdata_save	[	160	]	<=	tdata_save	[	160	]	;
					tdata_save	[	161	]	<=	tdata_save	[	161	]	;
					tdata_save	[	162	]	<=	tdata_save	[	162	]	;
					tdata_save	[	163	]	<=	tdata_save	[	163	]	;
					tdata_save	[	164	]	<=	tdata_save	[	164	]	;
					tdata_save	[	165	]	<=	tdata_save	[	165	]	;
					tdata_save	[	166	]	<=	tdata_save	[	166	]	;
					tdata_save	[	167	]	<=	tdata_save	[	167	]	;
					tdata_save	[	168	]	<=	tdata_save	[	168	]	;
					tdata_save	[	169	]	<=	tdata_save	[	169	]	;
					tdata_save	[	170	]	<=	tdata_save	[	170	]	;
					tdata_save	[	171	]	<=	tdata_save	[	171	]	;
					tdata_save	[	172	]	<=	tdata_save	[	172	]	;
					tdata_save	[	173	]	<=	tdata_save	[	173	]	;
					tdata_save	[	174	]	<=	tdata_save	[	174	]	;
					tdata_save	[	175	]	<=	tdata_save	[	175	]	;
					tdata_save	[	176	]	<=	tdata_save	[	176	]	;
					tdata_save	[	177	]	<=	tdata_save	[	177	]	;
					tdata_save	[	178	]	<=	tdata_save	[	178	]	;
					tdata_save	[	179	]	<=	tdata_save	[	179	]	;
					tdata_save	[	180	]	<=	tdata_save	[	180	]	;
					tdata_save	[	181	]	<=	tdata_save	[	181	]	;
					tdata_save	[	182	]	<=	tdata_save	[	182	]	;
					tdata_save	[	183	]	<=	tdata_save	[	183	]	;
					tdata_save	[	184	]	<=	tdata_save	[	184	]	;
					tdata_save	[	185	]	<=	tdata_save	[	185	]	;
					tdata_save	[	186	]	<=	tdata_save	[	186	]	;
					tdata_save	[	187	]	<=	tdata_save	[	187	]	;
					tdata_save	[	188	]	<=	tdata_save	[	188	]	;
					tdata_save	[	189	]	<=	tdata_save	[	189	]	;
					tdata_save	[	190	]	<=	tdata_save	[	190	]	;
					tdata_save	[	191	]	<=	tdata_save	[	191	]	;
					tdata_save	[	192	]	<=	tdata_save	[	192	]	;
					tdata_save	[	193	]	<=	tdata_save	[	193	]	;
					tdata_save	[	194	]	<=	tdata_save	[	194	]	;
					tdata_save	[	195	]	<=	tdata_save	[	195	]	;
					tdata_save	[	196	]	<=	tdata_save	[	196	]	;
					tdata_save	[	197	]	<=	tdata_save	[	197	]	;
					tdata_save	[	198	]	<=	tdata_save	[	198	]	;
					tdata_save	[	199	]	<=	tdata_save	[	199	]	;
					tdata_save	[	200	]	<=	tdata_save	[	200	]	;
					tdata_save	[	201	]	<=	tdata_save	[	201	]	;
					tdata_save	[	202	]	<=	tdata_save	[	202	]	;
					tdata_save	[	203	]	<=	tdata_save	[	203	]	;
					tdata_save	[	204	]	<=	tdata_save	[	204	]	;
					tdata_save	[	205	]	<=	tdata_save	[	205	]	;
					tdata_save	[	206	]	<=	tdata_save	[	206	]	;
					tdata_save	[	207	]	<=	tdata_save	[	207	]	;
					tdata_save	[	208	]	<=	tdata_save	[	208	]	;
					tdata_save	[	209	]	<=	tdata_save	[	209	]	;
					tdata_save	[	210	]	<=	tdata_save	[	210	]	;
					tdata_save	[	211	]	<=	tdata_save	[	211	]	;
					tdata_save	[	212	]	<=	tdata_save	[	212	]	;
					tdata_save	[	213	]	<=	tdata_save	[	213	]	;
					tdata_save	[	214	]	<=	tdata_save	[	214	]	;
					tdata_save	[	215	]	<=	tdata_save	[	215	]	;
					tdata_save	[	216	]	<=	tdata_save	[	216	]	;
					tdata_save	[	217	]	<=	tdata_save	[	217	]	;
					tdata_save	[	218	]	<=	tdata_save	[	218	]	;
					tdata_save	[	219	]	<=	tdata_save	[	219	]	;
					tdata_save	[	220	]	<=	tdata_save	[	220	]	;
					tdata_save	[	221	]	<=	tdata_save	[	221	]	;
					tdata_save	[	222	]	<=	tdata_save	[	222	]	;
					tdata_save	[	223	]	<=	tdata_save	[	223	]	;
					tdata_save	[	224	]	<=	tdata_save	[	224	]	;
					tdata_save	[	225	]	<=	tdata_save	[	225	]	;
					tdata_save	[	226	]	<=	tdata_save	[	226	]	;
					tdata_save	[	227	]	<=	tdata_save	[	227	]	;
					tdata_save	[	228	]	<=	tdata_save	[	228	]	;
					tdata_save	[	229	]	<=	tdata_save	[	229	]	;
					tdata_save	[	230	]	<=	tdata_save	[	230	]	;
					tdata_save	[	231	]	<=	tdata_save	[	231	]	;
					tdata_save	[	232	]	<=	tdata_save	[	232	]	;
					tdata_save	[	233	]	<=	tdata_save	[	233	]	;
					tdata_save	[	234	]	<=	tdata_save	[	234	]	;
					tdata_save	[	235	]	<=	tdata_save	[	235	]	;
					tdata_save	[	236	]	<=	tdata_save	[	236	]	;
					tdata_save	[	237	]	<=	tdata_save	[	237	]	;
					tdata_save	[	238	]	<=	tdata_save	[	238	]	;
					tdata_save	[	239	]	<=	tdata_save	[	239	]	;
					tdata_save	[	240	]	<=	tdata_save	[	240	]	;
					tdata_save	[	241	]	<=	tdata_save	[	241	]	;
					tdata_save	[	242	]	<=	tdata_save	[	242	]	;
					tdata_save	[	243	]	<=	tdata_save	[	243	]	;
					tdata_save	[	244	]	<=	tdata_save	[	244	]	;
					tdata_save	[	245	]	<=	tdata_save	[	245	]	;
					tdata_save	[	246	]	<=	tdata_save	[	246	]	;
					tdata_save	[	247	]	<=	tdata_save	[	247	]	;
					tdata_save	[	248	]	<=	tdata_save	[	248	]	;
					tdata_save	[	249	]	<=	tdata_save	[	249	]	;
					tdata_save	[	250	]	<=	tdata_save	[	250	]	;
					tdata_save	[	251	]	<=	tdata_save	[	251	]	;
					tdata_save	[	252	]	<=	tdata_save	[	252	]	;
					tdata_save	[	253	]	<=	tdata_save	[	253	]	;
					tdata_save	[	254	]	<=	tdata_save	[	254	]	;
					tdata_save	[	255	]	<=	tdata_save	[	255	]	;
									tuser_save	[	0	]	<=	tuser_save	[	0	]	;
				tuser_save	[	1	]	<=	tuser_save	[	1	]	;
				tuser_save	[	2	]	<=	tuser_save	[	2	]	;
				tuser_save	[	3	]	<=	tuser_save	[	3	]	;
				tuser_save	[	4	]	<=	tuser_save	[	4	]	;
				tuser_save	[	5	]	<=	tuser_save	[	5	]	;
				tuser_save	[	6	]	<=	tuser_save	[	6	]	;
				tuser_save	[	7	]	<=	tuser_save	[	7	]	;
				tuser_save	[	8	]	<=	tuser_save	[	8	]	;
				tuser_save	[	9	]	<=	tuser_save	[	9	]	;
				tuser_save	[	10	]	<=	tuser_save	[	10	]	;
				tuser_save	[	11	]	<=	tuser_save	[	11	]	;
				tuser_save	[	12	]	<=	tuser_save	[	12	]	;
				tuser_save	[	13	]	<=	tuser_save	[	13	]	;
				tuser_save	[	14	]	<=	tuser_save	[	14	]	;
				tuser_save	[	15	]	<=	tuser_save	[	15	]	;
				tuser_save	[	16	]	<=	tuser_save	[	16	]	;
				tuser_save	[	17	]	<=	tuser_save	[	17	]	;
				tuser_save	[	18	]	<=	tuser_save	[	18	]	;
				tuser_save	[	19	]	<=	tuser_save	[	19	]	;
				tuser_save	[	20	]	<=	tuser_save	[	20	]	;
				tuser_save	[	21	]	<=	tuser_save	[	21	]	;
				tuser_save	[	22	]	<=	tuser_save	[	22	]	;
				tuser_save	[	23	]	<=	tuser_save	[	23	]	;
				tuser_save	[	24	]	<=	tuser_save	[	24	]	;
				tuser_save	[	25	]	<=	tuser_save	[	25	]	;
				tuser_save	[	26	]	<=	tuser_save	[	26	]	;
				tuser_save	[	27	]	<=	tuser_save	[	27	]	;
				tuser_save	[	28	]	<=	tuser_save	[	28	]	;
				tuser_save	[	29	]	<=	tuser_save	[	29	]	;
				tuser_save	[	30	]	<=	tuser_save	[	30	]	;
				tuser_save	[	31	]	<=	tuser_save	[	31	]	;
				tuser_save	[	32	]	<=	tuser_save	[	32	]	;
				tuser_save	[	33	]	<=	tuser_save	[	33	]	;
				tuser_save	[	34	]	<=	tuser_save	[	34	]	;
				tuser_save	[	35	]	<=	tuser_save	[	35	]	;
				tuser_save	[	36	]	<=	tuser_save	[	36	]	;
				tuser_save	[	37	]	<=	tuser_save	[	37	]	;
				tuser_save	[	38	]	<=	tuser_save	[	38	]	;
				tuser_save	[	39	]	<=	tuser_save	[	39	]	;
				tuser_save	[	40	]	<=	tuser_save	[	40	]	;
				tuser_save	[	41	]	<=	tuser_save	[	41	]	;
				tuser_save	[	42	]	<=	tuser_save	[	42	]	;
				tuser_save	[	43	]	<=	tuser_save	[	43	]	;
				tuser_save	[	44	]	<=	tuser_save	[	44	]	;
				tuser_save	[	45	]	<=	tuser_save	[	45	]	;
				tuser_save	[	46	]	<=	tuser_save	[	46	]	;
				tuser_save	[	47	]	<=	tuser_save	[	47	]	;
				tuser_save	[	48	]	<=	tuser_save	[	48	]	;
				tuser_save	[	49	]	<=	tuser_save	[	49	]	;
				tuser_save	[	50	]	<=	tuser_save	[	50	]	;
				tuser_save	[	51	]	<=	tuser_save	[	51	]	;
				tuser_save	[	52	]	<=	tuser_save	[	52	]	;
				tuser_save	[	53	]	<=	tuser_save	[	53	]	;
				tuser_save	[	54	]	<=	tuser_save	[	54	]	;
				tuser_save	[	55	]	<=	tuser_save	[	55	]	;
				tuser_save	[	56	]	<=	tuser_save	[	56	]	;
				tuser_save	[	57	]	<=	tuser_save	[	57	]	;
				tuser_save	[	58	]	<=	tuser_save	[	58	]	;
				tuser_save	[	59	]	<=	tuser_save	[	59	]	;
				tuser_save	[	60	]	<=	tuser_save	[	60	]	;
				tuser_save	[	61	]	<=	tuser_save	[	61	]	;
				tuser_save	[	62	]	<=	tuser_save	[	62	]	;
				tuser_save	[	63	]	<=	tuser_save	[	63	]	;
				tuser_save	[	64	]	<=	tuser_save	[	64	]	;
				tuser_save	[	65	]	<=	tuser_save	[	65	]	;
				tuser_save	[	66	]	<=	tuser_save	[	66	]	;
				tuser_save	[	67	]	<=	tuser_save	[	67	]	;
				tuser_save	[	68	]	<=	tuser_save	[	68	]	;
				tuser_save	[	69	]	<=	tuser_save	[	69	]	;
				tuser_save	[	70	]	<=	tuser_save	[	70	]	;
				tuser_save	[	71	]	<=	tuser_save	[	71	]	;
				tuser_save	[	72	]	<=	tuser_save	[	72	]	;
				tuser_save	[	73	]	<=	tuser_save	[	73	]	;
				tuser_save	[	74	]	<=	tuser_save	[	74	]	;
				tuser_save	[	75	]	<=	tuser_save	[	75	]	;
				tuser_save	[	76	]	<=	tuser_save	[	76	]	;
				tuser_save	[	77	]	<=	tuser_save	[	77	]	;
				tuser_save	[	78	]	<=	tuser_save	[	78	]	;
				tuser_save	[	79	]	<=	tuser_save	[	79	]	;
				tuser_save	[	80	]	<=	tuser_save	[	80	]	;
				tuser_save	[	81	]	<=	tuser_save	[	81	]	;
				tuser_save	[	82	]	<=	tuser_save	[	82	]	;
				tuser_save	[	83	]	<=	tuser_save	[	83	]	;
				tuser_save	[	84	]	<=	tuser_save	[	84	]	;
				tuser_save	[	85	]	<=	tuser_save	[	85	]	;
				tuser_save	[	86	]	<=	tuser_save	[	86	]	;
				tuser_save	[	87	]	<=	tuser_save	[	87	]	;
				tuser_save	[	88	]	<=	tuser_save	[	88	]	;
				tuser_save	[	89	]	<=	tuser_save	[	89	]	;
				tuser_save	[	90	]	<=	tuser_save	[	90	]	;
				tuser_save	[	91	]	<=	tuser_save	[	91	]	;
				tuser_save	[	92	]	<=	tuser_save	[	92	]	;
				tuser_save	[	93	]	<=	tuser_save	[	93	]	;
				tuser_save	[	94	]	<=	tuser_save	[	94	]	;
				tuser_save	[	95	]	<=	tuser_save	[	95	]	;
				tuser_save	[	96	]	<=	tuser_save	[	96	]	;
				tuser_save	[	97	]	<=	tuser_save	[	97	]	;
				tuser_save	[	98	]	<=	tuser_save	[	98	]	;
				tuser_save	[	99	]	<=	tuser_save	[	99	]	;
				tuser_save	[	100	]	<=	tuser_save	[	100	]	;
				tuser_save	[	101	]	<=	tuser_save	[	101	]	;
				tuser_save	[	102	]	<=	tuser_save	[	102	]	;
				tuser_save	[	103	]	<=	tuser_save	[	103	]	;
				tuser_save	[	104	]	<=	tuser_save	[	104	]	;
				tuser_save	[	105	]	<=	tuser_save	[	105	]	;
				tuser_save	[	106	]	<=	tuser_save	[	106	]	;
				tuser_save	[	107	]	<=	tuser_save	[	107	]	;
				tuser_save	[	108	]	<=	tuser_save	[	108	]	;
				tuser_save	[	109	]	<=	tuser_save	[	109	]	;
				tuser_save	[	110	]	<=	tuser_save	[	110	]	;
				tuser_save	[	111	]	<=	tuser_save	[	111	]	;
				tuser_save	[	112	]	<=	tuser_save	[	112	]	;
				tuser_save	[	113	]	<=	tuser_save	[	113	]	;
				tuser_save	[	114	]	<=	tuser_save	[	114	]	;
				tuser_save	[	115	]	<=	tuser_save	[	115	]	;
				tuser_save	[	116	]	<=	tuser_save	[	116	]	;
				tuser_save	[	117	]	<=	tuser_save	[	117	]	;
				tuser_save	[	118	]	<=	tuser_save	[	118	]	;
				tuser_save	[	119	]	<=	tuser_save	[	119	]	;
				tuser_save	[	120	]	<=	tuser_save	[	120	]	;
				tuser_save	[	121	]	<=	tuser_save	[	121	]	;
				tuser_save	[	122	]	<=	tuser_save	[	122	]	;
				tuser_save	[	123	]	<=	tuser_save	[	123	]	;
				tuser_save	[	124	]	<=	tuser_save	[	124	]	;
				tuser_save	[	125	]	<=	tuser_save	[	125	]	;
				tuser_save	[	126	]	<=	tuser_save	[	126	]	;
				tuser_save	[	127	]	<=	tuser_save	[	127	]	;
				tuser_save	[	128	]	<=	tuser_save	[	128	]	;
				tuser_save	[	129	]	<=	tuser_save	[	129	]	;
				tuser_save	[	130	]	<=	tuser_save	[	130	]	;
				tuser_save	[	131	]	<=	tuser_save	[	131	]	;
				tuser_save	[	132	]	<=	tuser_save	[	132	]	;
				tuser_save	[	133	]	<=	tuser_save	[	133	]	;
				tuser_save	[	134	]	<=	tuser_save	[	134	]	;
				tuser_save	[	135	]	<=	tuser_save	[	135	]	;
				tuser_save	[	136	]	<=	tuser_save	[	136	]	;
				tuser_save	[	137	]	<=	tuser_save	[	137	]	;
				tuser_save	[	138	]	<=	tuser_save	[	138	]	;
				tuser_save	[	139	]	<=	tuser_save	[	139	]	;
				tuser_save	[	140	]	<=	tuser_save	[	140	]	;
				tuser_save	[	141	]	<=	tuser_save	[	141	]	;
				tuser_save	[	142	]	<=	tuser_save	[	142	]	;
				tuser_save	[	143	]	<=	tuser_save	[	143	]	;
				tuser_save	[	144	]	<=	tuser_save	[	144	]	;
				tuser_save	[	145	]	<=	tuser_save	[	145	]	;
				tuser_save	[	146	]	<=	tuser_save	[	146	]	;
				tuser_save	[	147	]	<=	tuser_save	[	147	]	;
				tuser_save	[	148	]	<=	tuser_save	[	148	]	;
				tuser_save	[	149	]	<=	tuser_save	[	149	]	;
				tuser_save	[	150	]	<=	tuser_save	[	150	]	;
				tuser_save	[	151	]	<=	tuser_save	[	151	]	;
				tuser_save	[	152	]	<=	tuser_save	[	152	]	;
				tuser_save	[	153	]	<=	tuser_save	[	153	]	;
				tuser_save	[	154	]	<=	tuser_save	[	154	]	;
				tuser_save	[	155	]	<=	tuser_save	[	155	]	;
				tuser_save	[	156	]	<=	tuser_save	[	156	]	;
				tuser_save	[	157	]	<=	tuser_save	[	157	]	;
				tuser_save	[	158	]	<=	tuser_save	[	158	]	;
				tuser_save	[	159	]	<=	tuser_save	[	159	]	;
				tuser_save	[	160	]	<=	tuser_save	[	160	]	;
				tuser_save	[	161	]	<=	tuser_save	[	161	]	;
				tuser_save	[	162	]	<=	tuser_save	[	162	]	;
				tuser_save	[	163	]	<=	tuser_save	[	163	]	;
				tuser_save	[	164	]	<=	tuser_save	[	164	]	;
				tuser_save	[	165	]	<=	tuser_save	[	165	]	;
				tuser_save	[	166	]	<=	tuser_save	[	166	]	;
				tuser_save	[	167	]	<=	tuser_save	[	167	]	;
				tuser_save	[	168	]	<=	tuser_save	[	168	]	;
				tuser_save	[	169	]	<=	tuser_save	[	169	]	;
				tuser_save	[	170	]	<=	tuser_save	[	170	]	;
				tuser_save	[	171	]	<=	tuser_save	[	171	]	;
				tuser_save	[	172	]	<=	tuser_save	[	172	]	;
				tuser_save	[	173	]	<=	tuser_save	[	173	]	;
				tuser_save	[	174	]	<=	tuser_save	[	174	]	;
				tuser_save	[	175	]	<=	tuser_save	[	175	]	;
				tuser_save	[	176	]	<=	tuser_save	[	176	]	;
				tuser_save	[	177	]	<=	tuser_save	[	177	]	;
				tuser_save	[	178	]	<=	tuser_save	[	178	]	;
				tuser_save	[	179	]	<=	tuser_save	[	179	]	;
				tuser_save	[	180	]	<=	tuser_save	[	180	]	;
				tuser_save	[	181	]	<=	tuser_save	[	181	]	;
				tuser_save	[	182	]	<=	tuser_save	[	182	]	;
				tuser_save	[	183	]	<=	tuser_save	[	183	]	;
				tuser_save	[	184	]	<=	tuser_save	[	184	]	;
				tuser_save	[	185	]	<=	tuser_save	[	185	]	;
				tuser_save	[	186	]	<=	tuser_save	[	186	]	;
				tuser_save	[	187	]	<=	tuser_save	[	187	]	;
				tuser_save	[	188	]	<=	tuser_save	[	188	]	;
				tuser_save	[	189	]	<=	tuser_save	[	189	]	;
				tuser_save	[	190	]	<=	tuser_save	[	190	]	;
				tuser_save	[	191	]	<=	tuser_save	[	191	]	;
				tuser_save	[	192	]	<=	tuser_save	[	192	]	;
				tuser_save	[	193	]	<=	tuser_save	[	193	]	;
				tuser_save	[	194	]	<=	tuser_save	[	194	]	;
				tuser_save	[	195	]	<=	tuser_save	[	195	]	;
				tuser_save	[	196	]	<=	tuser_save	[	196	]	;
				tuser_save	[	197	]	<=	tuser_save	[	197	]	;
				tuser_save	[	198	]	<=	tuser_save	[	198	]	;
				tuser_save	[	199	]	<=	tuser_save	[	199	]	;
				tuser_save	[	200	]	<=	tuser_save	[	200	]	;
				tuser_save	[	201	]	<=	tuser_save	[	201	]	;
				tuser_save	[	202	]	<=	tuser_save	[	202	]	;
				tuser_save	[	203	]	<=	tuser_save	[	203	]	;
				tuser_save	[	204	]	<=	tuser_save	[	204	]	;
				tuser_save	[	205	]	<=	tuser_save	[	205	]	;
				tuser_save	[	206	]	<=	tuser_save	[	206	]	;
				tuser_save	[	207	]	<=	tuser_save	[	207	]	;
				tuser_save	[	208	]	<=	tuser_save	[	208	]	;
				tuser_save	[	209	]	<=	tuser_save	[	209	]	;
				tuser_save	[	210	]	<=	tuser_save	[	210	]	;
				tuser_save	[	211	]	<=	tuser_save	[	211	]	;
				tuser_save	[	212	]	<=	tuser_save	[	212	]	;
				tuser_save	[	213	]	<=	tuser_save	[	213	]	;
				tuser_save	[	214	]	<=	tuser_save	[	214	]	;
				tuser_save	[	215	]	<=	tuser_save	[	215	]	;
				tuser_save	[	216	]	<=	tuser_save	[	216	]	;
				tuser_save	[	217	]	<=	tuser_save	[	217	]	;
				tuser_save	[	218	]	<=	tuser_save	[	218	]	;
				tuser_save	[	219	]	<=	tuser_save	[	219	]	;
				tuser_save	[	220	]	<=	tuser_save	[	220	]	;
				tuser_save	[	221	]	<=	tuser_save	[	221	]	;
				tuser_save	[	222	]	<=	tuser_save	[	222	]	;
				tuser_save	[	223	]	<=	tuser_save	[	223	]	;
				tuser_save	[	224	]	<=	tuser_save	[	224	]	;
				tuser_save	[	225	]	<=	tuser_save	[	225	]	;
				tuser_save	[	226	]	<=	tuser_save	[	226	]	;
				tuser_save	[	227	]	<=	tuser_save	[	227	]	;
				tuser_save	[	228	]	<=	tuser_save	[	228	]	;
				tuser_save	[	229	]	<=	tuser_save	[	229	]	;
				tuser_save	[	230	]	<=	tuser_save	[	230	]	;
				tuser_save	[	231	]	<=	tuser_save	[	231	]	;
				tuser_save	[	232	]	<=	tuser_save	[	232	]	;
				tuser_save	[	233	]	<=	tuser_save	[	233	]	;
				tuser_save	[	234	]	<=	tuser_save	[	234	]	;
				tuser_save	[	235	]	<=	tuser_save	[	235	]	;
				tuser_save	[	236	]	<=	tuser_save	[	236	]	;
				tuser_save	[	237	]	<=	tuser_save	[	237	]	;
				tuser_save	[	238	]	<=	tuser_save	[	238	]	;
				tuser_save	[	239	]	<=	tuser_save	[	239	]	;
				tuser_save	[	240	]	<=	tuser_save	[	240	]	;
				tuser_save	[	241	]	<=	tuser_save	[	241	]	;
				tuser_save	[	242	]	<=	tuser_save	[	242	]	;
				tuser_save	[	243	]	<=	tuser_save	[	243	]	;
				tuser_save	[	244	]	<=	tuser_save	[	244	]	;
				tuser_save	[	245	]	<=	tuser_save	[	245	]	;
				tuser_save	[	246	]	<=	tuser_save	[	246	]	;
				tuser_save	[	247	]	<=	tuser_save	[	247	]	;
				tuser_save	[	248	]	<=	tuser_save	[	248	]	;
				tuser_save	[	249	]	<=	tuser_save	[	249	]	;
				tuser_save	[	250	]	<=	tuser_save	[	250	]	;
				tuser_save	[	251	]	<=	tuser_save	[	251	]	;
				tuser_save	[	252	]	<=	tuser_save	[	252	]	;
				tuser_save	[	253	]	<=	tuser_save	[	253	]	;
				tuser_save	[	254	]	<=	tuser_save	[	254	]	;
				tuser_save	[	255	]	<=	tuser_save	[	255	]	;
					if(count_packet == 2'd2)
					begin
						count_packet <= 2'd0;
					end
					else
					begin
						count_packet	<= count_packet;
					end
					sum_tdata		<=	201'd0;
					sum_tuser		<=	128'd0;
					sum_tdata_valid		<=	1'b0;
					sum_tuser_valid		<=	1'b0;
				end
			end
			else
			begin
				if((eth_type == 16'h0800) && (count_packet == 2'd0))
				begin
					tdata_save	[	0	]	<=	axififo_din;	//shift			
					tdata_save	[	1	]	<=	tdata_save	[	0	]	;
					tdata_save	[	2	]	<=	tdata_save	[	1	]	;
					tdata_save	[	3	]	<=	tdata_save	[	2	]	;
					tdata_save	[	4	]	<=	tdata_save	[	3	]	;
					tdata_save	[	5	]	<=	tdata_save	[	4	]	;
					tdata_save	[	6	]	<=	tdata_save	[	5	]	;
					tdata_save	[	7	]	<=	tdata_save	[	6	]	;
					tdata_save	[	8	]	<=	tdata_save	[	7	]	;
					tdata_save	[	9	]	<=	tdata_save	[	8	]	;
					tdata_save	[	10	]	<=	tdata_save	[	9	]	;
					tdata_save	[	11	]	<=	tdata_save	[	10	]	;
					tdata_save	[	12	]	<=	tdata_save	[	11	]	;
					tdata_save	[	13	]	<=	tdata_save	[	12	]	;
					tdata_save	[	14	]	<=	tdata_save	[	13	]	;
					tdata_save	[	15	]	<=	tdata_save	[	14	]	;
					tdata_save	[	16	]	<=	tdata_save	[	15	]	;
					tdata_save	[	17	]	<=	tdata_save	[	16	]	;
					tdata_save	[	18	]	<=	tdata_save	[	17	]	;
					tdata_save	[	19	]	<=	tdata_save	[	18	]	;
					tdata_save	[	20	]	<=	tdata_save	[	19	]	;
					tdata_save	[	21	]	<=	tdata_save	[	20	]	;
					tdata_save	[	22	]	<=	tdata_save	[	21	]	;
					tdata_save	[	23	]	<=	tdata_save	[	22	]	;
					tdata_save	[	24	]	<=	tdata_save	[	23	]	;
					tdata_save	[	25	]	<=	tdata_save	[	24	]	;
					tdata_save	[	26	]	<=	tdata_save	[	25	]	;
					tdata_save	[	27	]	<=	tdata_save	[	26	]	;
					tdata_save	[	28	]	<=	tdata_save	[	27	]	;
					tdata_save	[	29	]	<=	tdata_save	[	28	]	;
					tdata_save	[	30	]	<=	tdata_save	[	29	]	;
					tdata_save	[	31	]	<=	tdata_save	[	30	]	;
					tdata_save	[	32	]	<=	tdata_save	[	31	]	;
					tdata_save	[	33	]	<=	tdata_save	[	32	]	;
					tdata_save	[	34	]	<=	tdata_save	[	33	]	;
					tdata_save	[	35	]	<=	tdata_save	[	34	]	;
					tdata_save	[	36	]	<=	tdata_save	[	35	]	;
					tdata_save	[	37	]	<=	tdata_save	[	36	]	;
					tdata_save	[	38	]	<=	tdata_save	[	37	]	;
					tdata_save	[	39	]	<=	tdata_save	[	38	]	;
					tdata_save	[	40	]	<=	tdata_save	[	39	]	;
					tdata_save	[	41	]	<=	tdata_save	[	40	]	;
					tdata_save	[	42	]	<=	tdata_save	[	41	]	;
					tdata_save	[	43	]	<=	tdata_save	[	42	]	;
					tdata_save	[	44	]	<=	tdata_save	[	43	]	;
					tdata_save	[	45	]	<=	tdata_save	[	44	]	;
					tdata_save	[	46	]	<=	tdata_save	[	45	]	;
					tdata_save	[	47	]	<=	tdata_save	[	46	]	;
					tdata_save	[	48	]	<=	tdata_save	[	47	]	;
					tdata_save	[	49	]	<=	tdata_save	[	48	]	;
					tdata_save	[	50	]	<=	tdata_save	[	49	]	;
					tdata_save	[	51	]	<=	tdata_save	[	50	]	;
					tdata_save	[	52	]	<=	tdata_save	[	51	]	;
					tdata_save	[	53	]	<=	tdata_save	[	52	]	;
					tdata_save	[	54	]	<=	tdata_save	[	53	]	;
					tdata_save	[	55	]	<=	tdata_save	[	54	]	;
					tdata_save	[	56	]	<=	tdata_save	[	55	]	;
					tdata_save	[	57	]	<=	tdata_save	[	56	]	;
					tdata_save	[	58	]	<=	tdata_save	[	57	]	;
					tdata_save	[	59	]	<=	tdata_save	[	58	]	;
					tdata_save	[	60	]	<=	tdata_save	[	59	]	;
					tdata_save	[	61	]	<=	tdata_save	[	60	]	;
					tdata_save	[	62	]	<=	tdata_save	[	61	]	;
					tdata_save	[	63	]	<=	tdata_save	[	62	]	;
					tdata_save	[	64	]	<=	tdata_save	[	63	]	;
					tdata_save	[	65	]	<=	tdata_save	[	64	]	;
					tdata_save	[	66	]	<=	tdata_save	[	65	]	;
					tdata_save	[	67	]	<=	tdata_save	[	66	]	;
					tdata_save	[	68	]	<=	tdata_save	[	67	]	;
					tdata_save	[	69	]	<=	tdata_save	[	68	]	;
					tdata_save	[	70	]	<=	tdata_save	[	69	]	;
					tdata_save	[	71	]	<=	tdata_save	[	70	]	;
					tdata_save	[	72	]	<=	tdata_save	[	71	]	;
					tdata_save	[	73	]	<=	tdata_save	[	72	]	;
					tdata_save	[	74	]	<=	tdata_save	[	73	]	;
					tdata_save	[	75	]	<=	tdata_save	[	74	]	;
					tdata_save	[	76	]	<=	tdata_save	[	75	]	;
					tdata_save	[	77	]	<=	tdata_save	[	76	]	;
					tdata_save	[	78	]	<=	tdata_save	[	77	]	;
					tdata_save	[	79	]	<=	tdata_save	[	78	]	;
					tdata_save	[	80	]	<=	tdata_save	[	79	]	;
					tdata_save	[	81	]	<=	tdata_save	[	80	]	;
					tdata_save	[	82	]	<=	tdata_save	[	81	]	;
					tdata_save	[	83	]	<=	tdata_save	[	82	]	;
					tdata_save	[	84	]	<=	tdata_save	[	83	]	;
					tdata_save	[	85	]	<=	tdata_save	[	84	]	;
					tdata_save	[	86	]	<=	tdata_save	[	85	]	;
					tdata_save	[	87	]	<=	tdata_save	[	86	]	;
					tdata_save	[	88	]	<=	tdata_save	[	87	]	;
					tdata_save	[	89	]	<=	tdata_save	[	88	]	;
					tdata_save	[	90	]	<=	tdata_save	[	89	]	;
					tdata_save	[	91	]	<=	tdata_save	[	90	]	;
					tdata_save	[	92	]	<=	tdata_save	[	91	]	;
					tdata_save	[	93	]	<=	tdata_save	[	92	]	;
					tdata_save	[	94	]	<=	tdata_save	[	93	]	;
					tdata_save	[	95	]	<=	tdata_save	[	94	]	;
					tdata_save	[	96	]	<=	tdata_save	[	95	]	;
					tdata_save	[	97	]	<=	tdata_save	[	96	]	;
					tdata_save	[	98	]	<=	tdata_save	[	97	]	;
					tdata_save	[	99	]	<=	tdata_save	[	98	]	;
					tdata_save	[	100	]	<=	tdata_save	[	99	]	;
					tdata_save	[	101	]	<=	tdata_save	[	100	]	;
					tdata_save	[	102	]	<=	tdata_save	[	101	]	;
					tdata_save	[	103	]	<=	tdata_save	[	102	]	;
					tdata_save	[	104	]	<=	tdata_save	[	103	]	;
					tdata_save	[	105	]	<=	tdata_save	[	104	]	;
					tdata_save	[	106	]	<=	tdata_save	[	105	]	;
					tdata_save	[	107	]	<=	tdata_save	[	106	]	;
					tdata_save	[	108	]	<=	tdata_save	[	107	]	;
					tdata_save	[	109	]	<=	tdata_save	[	108	]	;
					tdata_save	[	110	]	<=	tdata_save	[	109	]	;
					tdata_save	[	111	]	<=	tdata_save	[	110	]	;
					tdata_save	[	112	]	<=	tdata_save	[	111	]	;
					tdata_save	[	113	]	<=	tdata_save	[	112	]	;
					tdata_save	[	114	]	<=	tdata_save	[	113	]	;
					tdata_save	[	115	]	<=	tdata_save	[	114	]	;
					tdata_save	[	116	]	<=	tdata_save	[	115	]	;
					tdata_save	[	117	]	<=	tdata_save	[	116	]	;
					tdata_save	[	118	]	<=	tdata_save	[	117	]	;
					tdata_save	[	119	]	<=	tdata_save	[	118	]	;
					tdata_save	[	120	]	<=	tdata_save	[	119	]	;
					tdata_save	[	121	]	<=	tdata_save	[	120	]	;
					tdata_save	[	122	]	<=	tdata_save	[	121	]	;
					tdata_save	[	123	]	<=	tdata_save	[	122	]	;
					tdata_save	[	124	]	<=	tdata_save	[	123	]	;
					tdata_save	[	125	]	<=	tdata_save	[	124	]	;
					tdata_save	[	126	]	<=	tdata_save	[	125	]	;
					tdata_save	[	127	]	<=	tdata_save	[	126	]	;
					tdata_save	[	128	]	<=	tdata_save	[	127	]	;
					tdata_save	[	129	]	<=	tdata_save	[	128	]	;
					tdata_save	[	130	]	<=	tdata_save	[	129	]	;
					tdata_save	[	131	]	<=	tdata_save	[	130	]	;
					tdata_save	[	132	]	<=	tdata_save	[	131	]	;
					tdata_save	[	133	]	<=	tdata_save	[	132	]	;
					tdata_save	[	134	]	<=	tdata_save	[	133	]	;
					tdata_save	[	135	]	<=	tdata_save	[	134	]	;
					tdata_save	[	136	]	<=	tdata_save	[	135	]	;
					tdata_save	[	137	]	<=	tdata_save	[	136	]	;
					tdata_save	[	138	]	<=	tdata_save	[	137	]	;
					tdata_save	[	139	]	<=	tdata_save	[	138	]	;
					tdata_save	[	140	]	<=	tdata_save	[	139	]	;
					tdata_save	[	141	]	<=	tdata_save	[	140	]	;
					tdata_save	[	142	]	<=	tdata_save	[	141	]	;
					tdata_save	[	143	]	<=	tdata_save	[	142	]	;
					tdata_save	[	144	]	<=	tdata_save	[	143	]	;
					tdata_save	[	145	]	<=	tdata_save	[	144	]	;
					tdata_save	[	146	]	<=	tdata_save	[	145	]	;
					tdata_save	[	147	]	<=	tdata_save	[	146	]	;
					tdata_save	[	148	]	<=	tdata_save	[	147	]	;
					tdata_save	[	149	]	<=	tdata_save	[	148	]	;
					tdata_save	[	150	]	<=	tdata_save	[	149	]	;
					tdata_save	[	151	]	<=	tdata_save	[	150	]	;
					tdata_save	[	152	]	<=	tdata_save	[	151	]	;
					tdata_save	[	153	]	<=	tdata_save	[	152	]	;
					tdata_save	[	154	]	<=	tdata_save	[	153	]	;
					tdata_save	[	155	]	<=	tdata_save	[	154	]	;
					tdata_save	[	156	]	<=	tdata_save	[	155	]	;
					tdata_save	[	157	]	<=	tdata_save	[	156	]	;
					tdata_save	[	158	]	<=	tdata_save	[	157	]	;
					tdata_save	[	159	]	<=	tdata_save	[	158	]	;
					tdata_save	[	160	]	<=	tdata_save	[	159	]	;
					tdata_save	[	161	]	<=	tdata_save	[	160	]	;
					tdata_save	[	162	]	<=	tdata_save	[	161	]	;
					tdata_save	[	163	]	<=	tdata_save	[	162	]	;
					tdata_save	[	164	]	<=	tdata_save	[	163	]	;
					tdata_save	[	165	]	<=	tdata_save	[	164	]	;
					tdata_save	[	166	]	<=	tdata_save	[	165	]	;
					tdata_save	[	167	]	<=	tdata_save	[	166	]	;
					tdata_save	[	168	]	<=	tdata_save	[	167	]	;
					tdata_save	[	169	]	<=	tdata_save	[	168	]	;
					tdata_save	[	170	]	<=	tdata_save	[	169	]	;
					tdata_save	[	171	]	<=	tdata_save	[	170	]	;
					tdata_save	[	172	]	<=	tdata_save	[	171	]	;
					tdata_save	[	173	]	<=	tdata_save	[	172	]	;
					tdata_save	[	174	]	<=	tdata_save	[	173	]	;
					tdata_save	[	175	]	<=	tdata_save	[	174	]	;
					tdata_save	[	176	]	<=	tdata_save	[	175	]	;
					tdata_save	[	177	]	<=	tdata_save	[	176	]	;
					tdata_save	[	178	]	<=	tdata_save	[	177	]	;
					tdata_save	[	179	]	<=	tdata_save	[	178	]	;
					tdata_save	[	180	]	<=	tdata_save	[	179	]	;
					tdata_save	[	181	]	<=	tdata_save	[	180	]	;
					tdata_save	[	182	]	<=	tdata_save	[	181	]	;
					tdata_save	[	183	]	<=	tdata_save	[	182	]	;
					tdata_save	[	184	]	<=	tdata_save	[	183	]	;
					tdata_save	[	185	]	<=	tdata_save	[	184	]	;
					tdata_save	[	186	]	<=	tdata_save	[	185	]	;
					tdata_save	[	187	]	<=	tdata_save	[	186	]	;
					tdata_save	[	188	]	<=	tdata_save	[	187	]	;
					tdata_save	[	189	]	<=	tdata_save	[	188	]	;
					tdata_save	[	190	]	<=	tdata_save	[	189	]	;
					tdata_save	[	191	]	<=	tdata_save	[	190	]	;
					tdata_save	[	192	]	<=	tdata_save	[	191	]	;
					tdata_save	[	193	]	<=	tdata_save	[	192	]	;
					tdata_save	[	194	]	<=	tdata_save	[	193	]	;
					tdata_save	[	195	]	<=	tdata_save	[	194	]	;
					tdata_save	[	196	]	<=	tdata_save	[	195	]	;
					tdata_save	[	197	]	<=	tdata_save	[	196	]	;
					tdata_save	[	198	]	<=	tdata_save	[	197	]	;
					tdata_save	[	199	]	<=	tdata_save	[	198	]	;
					tdata_save	[	200	]	<=	tdata_save	[	199	]	;
					tdata_save	[	201	]	<=	tdata_save	[	200	]	;
					tdata_save	[	202	]	<=	tdata_save	[	201	]	;
					tdata_save	[	203	]	<=	tdata_save	[	202	]	;
					tdata_save	[	204	]	<=	tdata_save	[	203	]	;
					tdata_save	[	205	]	<=	tdata_save	[	204	]	;
					tdata_save	[	206	]	<=	tdata_save	[	205	]	;
					tdata_save	[	207	]	<=	tdata_save	[	206	]	;
					tdata_save	[	208	]	<=	tdata_save	[	207	]	;
					tdata_save	[	209	]	<=	tdata_save	[	208	]	;
					tdata_save	[	210	]	<=	tdata_save	[	209	]	;
					tdata_save	[	211	]	<=	tdata_save	[	210	]	;
					tdata_save	[	212	]	<=	tdata_save	[	211	]	;
					tdata_save	[	213	]	<=	tdata_save	[	212	]	;
					tdata_save	[	214	]	<=	tdata_save	[	213	]	;
					tdata_save	[	215	]	<=	tdata_save	[	214	]	;
					tdata_save	[	216	]	<=	tdata_save	[	215	]	;
					tdata_save	[	217	]	<=	tdata_save	[	216	]	;
					tdata_save	[	218	]	<=	tdata_save	[	217	]	;
					tdata_save	[	219	]	<=	tdata_save	[	218	]	;
					tdata_save	[	220	]	<=	tdata_save	[	219	]	;
					tdata_save	[	221	]	<=	tdata_save	[	220	]	;
					tdata_save	[	222	]	<=	tdata_save	[	221	]	;
					tdata_save	[	223	]	<=	tdata_save	[	222	]	;
					tdata_save	[	224	]	<=	tdata_save	[	223	]	;
					tdata_save	[	225	]	<=	tdata_save	[	224	]	;
					tdata_save	[	226	]	<=	tdata_save	[	225	]	;
					tdata_save	[	227	]	<=	tdata_save	[	226	]	;
					tdata_save	[	228	]	<=	tdata_save	[	227	]	;
					tdata_save	[	229	]	<=	tdata_save	[	228	]	;
					tdata_save	[	230	]	<=	tdata_save	[	229	]	;
					tdata_save	[	231	]	<=	tdata_save	[	230	]	;
					tdata_save	[	232	]	<=	tdata_save	[	231	]	;
					tdata_save	[	233	]	<=	tdata_save	[	232	]	;
					tdata_save	[	234	]	<=	tdata_save	[	233	]	;
					tdata_save	[	235	]	<=	tdata_save	[	234	]	;
					tdata_save	[	236	]	<=	tdata_save	[	235	]	;
					tdata_save	[	237	]	<=	tdata_save	[	236	]	;
					tdata_save	[	238	]	<=	tdata_save	[	237	]	;
					tdata_save	[	239	]	<=	tdata_save	[	238	]	;
					tdata_save	[	240	]	<=	tdata_save	[	239	]	;
					tdata_save	[	241	]	<=	tdata_save	[	240	]	;
					tdata_save	[	242	]	<=	tdata_save	[	241	]	;
					tdata_save	[	243	]	<=	tdata_save	[	242	]	;
					tdata_save	[	244	]	<=	tdata_save	[	243	]	;
					tdata_save	[	245	]	<=	tdata_save	[	244	]	;
					tdata_save	[	246	]	<=	tdata_save	[	245	]	;
					tdata_save	[	247	]	<=	tdata_save	[	246	]	;
					tdata_save	[	248	]	<=	tdata_save	[	247	]	;
					tdata_save	[	249	]	<=	tdata_save	[	248	]	;
					tdata_save	[	250	]	<=	tdata_save	[	249	]	;
					tdata_save	[	251	]	<=	tdata_save	[	250	]	;
					tdata_save	[	252	]	<=	tdata_save	[	251	]	;
					tdata_save	[	253	]	<=	tdata_save	[	252	]	;
					tdata_save	[	254	]	<=	tdata_save	[	253	]	;
					tdata_save	[	255	]	<=	tdata_save	[	254	]	;
					tuser_save	[	0	]	<=	tuser;						
				tuser_save	[	1	]	<=	tuser_save	[	0	]	;
				tuser_save	[	2	]	<=	tuser_save	[	1	]	;
				tuser_save	[	3	]	<=	tuser_save	[	2	]	;
				tuser_save	[	4	]	<=	tuser_save	[	3	]	;
				tuser_save	[	5	]	<=	tuser_save	[	4	]	;
				tuser_save	[	6	]	<=	tuser_save	[	5	]	;
				tuser_save	[	7	]	<=	tuser_save	[	6	]	;
				tuser_save	[	8	]	<=	tuser_save	[	7	]	;
				tuser_save	[	9	]	<=	tuser_save	[	8	]	;
				tuser_save	[	10	]	<=	tuser_save	[	9	]	;
				tuser_save	[	11	]	<=	tuser_save	[	10	]	;
				tuser_save	[	12	]	<=	tuser_save	[	11	]	;
				tuser_save	[	13	]	<=	tuser_save	[	12	]	;
				tuser_save	[	14	]	<=	tuser_save	[	13	]	;
				tuser_save	[	15	]	<=	tuser_save	[	14	]	;
				tuser_save	[	16	]	<=	tuser_save	[	15	]	;
				tuser_save	[	17	]	<=	tuser_save	[	16	]	;
				tuser_save	[	18	]	<=	tuser_save	[	17	]	;
				tuser_save	[	19	]	<=	tuser_save	[	18	]	;
				tuser_save	[	20	]	<=	tuser_save	[	19	]	;
				tuser_save	[	21	]	<=	tuser_save	[	20	]	;
				tuser_save	[	22	]	<=	tuser_save	[	21	]	;
				tuser_save	[	23	]	<=	tuser_save	[	22	]	;
				tuser_save	[	24	]	<=	tuser_save	[	23	]	;
				tuser_save	[	25	]	<=	tuser_save	[	24	]	;
				tuser_save	[	26	]	<=	tuser_save	[	25	]	;
				tuser_save	[	27	]	<=	tuser_save	[	26	]	;
				tuser_save	[	28	]	<=	tuser_save	[	27	]	;
				tuser_save	[	29	]	<=	tuser_save	[	28	]	;
				tuser_save	[	30	]	<=	tuser_save	[	29	]	;
				tuser_save	[	31	]	<=	tuser_save	[	30	]	;
				tuser_save	[	32	]	<=	tuser_save	[	31	]	;
				tuser_save	[	33	]	<=	tuser_save	[	32	]	;
				tuser_save	[	34	]	<=	tuser_save	[	33	]	;
				tuser_save	[	35	]	<=	tuser_save	[	34	]	;
				tuser_save	[	36	]	<=	tuser_save	[	35	]	;
				tuser_save	[	37	]	<=	tuser_save	[	36	]	;
				tuser_save	[	38	]	<=	tuser_save	[	37	]	;
				tuser_save	[	39	]	<=	tuser_save	[	38	]	;
				tuser_save	[	40	]	<=	tuser_save	[	39	]	;
				tuser_save	[	41	]	<=	tuser_save	[	40	]	;
				tuser_save	[	42	]	<=	tuser_save	[	41	]	;
				tuser_save	[	43	]	<=	tuser_save	[	42	]	;
				tuser_save	[	44	]	<=	tuser_save	[	43	]	;
				tuser_save	[	45	]	<=	tuser_save	[	44	]	;
				tuser_save	[	46	]	<=	tuser_save	[	45	]	;
				tuser_save	[	47	]	<=	tuser_save	[	46	]	;
				tuser_save	[	48	]	<=	tuser_save	[	47	]	;
				tuser_save	[	49	]	<=	tuser_save	[	48	]	;
				tuser_save	[	50	]	<=	tuser_save	[	49	]	;
				tuser_save	[	51	]	<=	tuser_save	[	50	]	;
				tuser_save	[	52	]	<=	tuser_save	[	51	]	;
				tuser_save	[	53	]	<=	tuser_save	[	52	]	;
				tuser_save	[	54	]	<=	tuser_save	[	53	]	;
				tuser_save	[	55	]	<=	tuser_save	[	54	]	;
				tuser_save	[	56	]	<=	tuser_save	[	55	]	;
				tuser_save	[	57	]	<=	tuser_save	[	56	]	;
				tuser_save	[	58	]	<=	tuser_save	[	57	]	;
				tuser_save	[	59	]	<=	tuser_save	[	58	]	;
				tuser_save	[	60	]	<=	tuser_save	[	59	]	;
				tuser_save	[	61	]	<=	tuser_save	[	60	]	;
				tuser_save	[	62	]	<=	tuser_save	[	61	]	;
				tuser_save	[	63	]	<=	tuser_save	[	62	]	;
				tuser_save	[	64	]	<=	tuser_save	[	63	]	;
				tuser_save	[	65	]	<=	tuser_save	[	64	]	;
				tuser_save	[	66	]	<=	tuser_save	[	65	]	;
				tuser_save	[	67	]	<=	tuser_save	[	66	]	;
				tuser_save	[	68	]	<=	tuser_save	[	67	]	;
				tuser_save	[	69	]	<=	tuser_save	[	68	]	;
				tuser_save	[	70	]	<=	tuser_save	[	69	]	;
				tuser_save	[	71	]	<=	tuser_save	[	70	]	;
				tuser_save	[	72	]	<=	tuser_save	[	71	]	;
				tuser_save	[	73	]	<=	tuser_save	[	72	]	;
				tuser_save	[	74	]	<=	tuser_save	[	73	]	;
				tuser_save	[	75	]	<=	tuser_save	[	74	]	;
				tuser_save	[	76	]	<=	tuser_save	[	75	]	;
				tuser_save	[	77	]	<=	tuser_save	[	76	]	;
				tuser_save	[	78	]	<=	tuser_save	[	77	]	;
				tuser_save	[	79	]	<=	tuser_save	[	78	]	;
				tuser_save	[	80	]	<=	tuser_save	[	79	]	;
				tuser_save	[	81	]	<=	tuser_save	[	80	]	;
				tuser_save	[	82	]	<=	tuser_save	[	81	]	;
				tuser_save	[	83	]	<=	tuser_save	[	82	]	;
				tuser_save	[	84	]	<=	tuser_save	[	83	]	;
				tuser_save	[	85	]	<=	tuser_save	[	84	]	;
				tuser_save	[	86	]	<=	tuser_save	[	85	]	;
				tuser_save	[	87	]	<=	tuser_save	[	86	]	;
				tuser_save	[	88	]	<=	tuser_save	[	87	]	;
				tuser_save	[	89	]	<=	tuser_save	[	88	]	;
				tuser_save	[	90	]	<=	tuser_save	[	89	]	;
				tuser_save	[	91	]	<=	tuser_save	[	90	]	;
				tuser_save	[	92	]	<=	tuser_save	[	91	]	;
				tuser_save	[	93	]	<=	tuser_save	[	92	]	;
				tuser_save	[	94	]	<=	tuser_save	[	93	]	;
				tuser_save	[	95	]	<=	tuser_save	[	94	]	;
				tuser_save	[	96	]	<=	tuser_save	[	95	]	;
				tuser_save	[	97	]	<=	tuser_save	[	96	]	;
				tuser_save	[	98	]	<=	tuser_save	[	97	]	;
				tuser_save	[	99	]	<=	tuser_save	[	98	]	;
				tuser_save	[	100	]	<=	tuser_save	[	99	]	;
				tuser_save	[	101	]	<=	tuser_save	[	100	]	;
				tuser_save	[	102	]	<=	tuser_save	[	101	]	;
				tuser_save	[	103	]	<=	tuser_save	[	102	]	;
				tuser_save	[	104	]	<=	tuser_save	[	103	]	;
				tuser_save	[	105	]	<=	tuser_save	[	104	]	;
				tuser_save	[	106	]	<=	tuser_save	[	105	]	;
				tuser_save	[	107	]	<=	tuser_save	[	106	]	;
				tuser_save	[	108	]	<=	tuser_save	[	107	]	;
				tuser_save	[	109	]	<=	tuser_save	[	108	]	;
				tuser_save	[	110	]	<=	tuser_save	[	109	]	;
				tuser_save	[	111	]	<=	tuser_save	[	110	]	;
				tuser_save	[	112	]	<=	tuser_save	[	111	]	;
				tuser_save	[	113	]	<=	tuser_save	[	112	]	;
				tuser_save	[	114	]	<=	tuser_save	[	113	]	;
				tuser_save	[	115	]	<=	tuser_save	[	114	]	;
				tuser_save	[	116	]	<=	tuser_save	[	115	]	;
				tuser_save	[	117	]	<=	tuser_save	[	116	]	;
				tuser_save	[	118	]	<=	tuser_save	[	117	]	;
				tuser_save	[	119	]	<=	tuser_save	[	118	]	;
				tuser_save	[	120	]	<=	tuser_save	[	119	]	;
				tuser_save	[	121	]	<=	tuser_save	[	120	]	;
				tuser_save	[	122	]	<=	tuser_save	[	121	]	;
				tuser_save	[	123	]	<=	tuser_save	[	122	]	;
				tuser_save	[	124	]	<=	tuser_save	[	123	]	;
				tuser_save	[	125	]	<=	tuser_save	[	124	]	;
				tuser_save	[	126	]	<=	tuser_save	[	125	]	;
				tuser_save	[	127	]	<=	tuser_save	[	126	]	;
				tuser_save	[	128	]	<=	tuser_save	[	127	]	;
				tuser_save	[	129	]	<=	tuser_save	[	128	]	;
				tuser_save	[	130	]	<=	tuser_save	[	129	]	;
				tuser_save	[	131	]	<=	tuser_save	[	130	]	;
				tuser_save	[	132	]	<=	tuser_save	[	131	]	;
				tuser_save	[	133	]	<=	tuser_save	[	132	]	;
				tuser_save	[	134	]	<=	tuser_save	[	133	]	;
				tuser_save	[	135	]	<=	tuser_save	[	134	]	;
				tuser_save	[	136	]	<=	tuser_save	[	135	]	;
				tuser_save	[	137	]	<=	tuser_save	[	136	]	;
				tuser_save	[	138	]	<=	tuser_save	[	137	]	;
				tuser_save	[	139	]	<=	tuser_save	[	138	]	;
				tuser_save	[	140	]	<=	tuser_save	[	139	]	;
				tuser_save	[	141	]	<=	tuser_save	[	140	]	;
				tuser_save	[	142	]	<=	tuser_save	[	141	]	;
				tuser_save	[	143	]	<=	tuser_save	[	142	]	;
				tuser_save	[	144	]	<=	tuser_save	[	143	]	;
				tuser_save	[	145	]	<=	tuser_save	[	144	]	;
				tuser_save	[	146	]	<=	tuser_save	[	145	]	;
				tuser_save	[	147	]	<=	tuser_save	[	146	]	;
				tuser_save	[	148	]	<=	tuser_save	[	147	]	;
				tuser_save	[	149	]	<=	tuser_save	[	148	]	;
				tuser_save	[	150	]	<=	tuser_save	[	149	]	;
				tuser_save	[	151	]	<=	tuser_save	[	150	]	;
				tuser_save	[	152	]	<=	tuser_save	[	151	]	;
				tuser_save	[	153	]	<=	tuser_save	[	152	]	;
				tuser_save	[	154	]	<=	tuser_save	[	153	]	;
				tuser_save	[	155	]	<=	tuser_save	[	154	]	;
				tuser_save	[	156	]	<=	tuser_save	[	155	]	;
				tuser_save	[	157	]	<=	tuser_save	[	156	]	;
				tuser_save	[	158	]	<=	tuser_save	[	157	]	;
				tuser_save	[	159	]	<=	tuser_save	[	158	]	;
				tuser_save	[	160	]	<=	tuser_save	[	159	]	;
				tuser_save	[	161	]	<=	tuser_save	[	160	]	;
				tuser_save	[	162	]	<=	tuser_save	[	161	]	;
				tuser_save	[	163	]	<=	tuser_save	[	162	]	;
				tuser_save	[	164	]	<=	tuser_save	[	163	]	;
				tuser_save	[	165	]	<=	tuser_save	[	164	]	;
				tuser_save	[	166	]	<=	tuser_save	[	165	]	;
				tuser_save	[	167	]	<=	tuser_save	[	166	]	;
				tuser_save	[	168	]	<=	tuser_save	[	167	]	;
				tuser_save	[	169	]	<=	tuser_save	[	168	]	;
				tuser_save	[	170	]	<=	tuser_save	[	169	]	;
				tuser_save	[	171	]	<=	tuser_save	[	170	]	;
				tuser_save	[	172	]	<=	tuser_save	[	171	]	;
				tuser_save	[	173	]	<=	tuser_save	[	172	]	;
				tuser_save	[	174	]	<=	tuser_save	[	173	]	;
				tuser_save	[	175	]	<=	tuser_save	[	174	]	;
				tuser_save	[	176	]	<=	tuser_save	[	175	]	;
				tuser_save	[	177	]	<=	tuser_save	[	176	]	;
				tuser_save	[	178	]	<=	tuser_save	[	177	]	;
				tuser_save	[	179	]	<=	tuser_save	[	178	]	;
				tuser_save	[	180	]	<=	tuser_save	[	179	]	;
				tuser_save	[	181	]	<=	tuser_save	[	180	]	;
				tuser_save	[	182	]	<=	tuser_save	[	181	]	;
				tuser_save	[	183	]	<=	tuser_save	[	182	]	;
				tuser_save	[	184	]	<=	tuser_save	[	183	]	;
				tuser_save	[	185	]	<=	tuser_save	[	184	]	;
				tuser_save	[	186	]	<=	tuser_save	[	185	]	;
				tuser_save	[	187	]	<=	tuser_save	[	186	]	;
				tuser_save	[	188	]	<=	tuser_save	[	187	]	;
				tuser_save	[	189	]	<=	tuser_save	[	188	]	;
				tuser_save	[	190	]	<=	tuser_save	[	189	]	;
				tuser_save	[	191	]	<=	tuser_save	[	190	]	;
				tuser_save	[	192	]	<=	tuser_save	[	191	]	;
				tuser_save	[	193	]	<=	tuser_save	[	192	]	;
				tuser_save	[	194	]	<=	tuser_save	[	193	]	;
				tuser_save	[	195	]	<=	tuser_save	[	194	]	;
				tuser_save	[	196	]	<=	tuser_save	[	195	]	;
				tuser_save	[	197	]	<=	tuser_save	[	196	]	;
				tuser_save	[	198	]	<=	tuser_save	[	197	]	;
				tuser_save	[	199	]	<=	tuser_save	[	198	]	;
				tuser_save	[	200	]	<=	tuser_save	[	199	]	;
				tuser_save	[	201	]	<=	tuser_save	[	200	]	;
				tuser_save	[	202	]	<=	tuser_save	[	201	]	;
				tuser_save	[	203	]	<=	tuser_save	[	202	]	;
				tuser_save	[	204	]	<=	tuser_save	[	203	]	;
				tuser_save	[	205	]	<=	tuser_save	[	204	]	;
				tuser_save	[	206	]	<=	tuser_save	[	205	]	;
				tuser_save	[	207	]	<=	tuser_save	[	206	]	;
				tuser_save	[	208	]	<=	tuser_save	[	207	]	;
				tuser_save	[	209	]	<=	tuser_save	[	208	]	;
				tuser_save	[	210	]	<=	tuser_save	[	209	]	;
				tuser_save	[	211	]	<=	tuser_save	[	210	]	;
				tuser_save	[	212	]	<=	tuser_save	[	211	]	;
				tuser_save	[	213	]	<=	tuser_save	[	212	]	;
				tuser_save	[	214	]	<=	tuser_save	[	213	]	;
				tuser_save	[	215	]	<=	tuser_save	[	214	]	;
				tuser_save	[	216	]	<=	tuser_save	[	215	]	;
				tuser_save	[	217	]	<=	tuser_save	[	216	]	;
				tuser_save	[	218	]	<=	tuser_save	[	217	]	;
				tuser_save	[	219	]	<=	tuser_save	[	218	]	;
				tuser_save	[	220	]	<=	tuser_save	[	219	]	;
				tuser_save	[	221	]	<=	tuser_save	[	220	]	;
				tuser_save	[	222	]	<=	tuser_save	[	221	]	;
				tuser_save	[	223	]	<=	tuser_save	[	222	]	;
				tuser_save	[	224	]	<=	tuser_save	[	223	]	;
				tuser_save	[	225	]	<=	tuser_save	[	224	]	;
				tuser_save	[	226	]	<=	tuser_save	[	225	]	;
				tuser_save	[	227	]	<=	tuser_save	[	226	]	;
				tuser_save	[	228	]	<=	tuser_save	[	227	]	;
				tuser_save	[	229	]	<=	tuser_save	[	228	]	;
				tuser_save	[	230	]	<=	tuser_save	[	229	]	;
				tuser_save	[	231	]	<=	tuser_save	[	230	]	;
				tuser_save	[	232	]	<=	tuser_save	[	231	]	;
				tuser_save	[	233	]	<=	tuser_save	[	232	]	;
				tuser_save	[	234	]	<=	tuser_save	[	233	]	;
				tuser_save	[	235	]	<=	tuser_save	[	234	]	;
				tuser_save	[	236	]	<=	tuser_save	[	235	]	;
				tuser_save	[	237	]	<=	tuser_save	[	236	]	;
				tuser_save	[	238	]	<=	tuser_save	[	237	]	;
				tuser_save	[	239	]	<=	tuser_save	[	238	]	;
				tuser_save	[	240	]	<=	tuser_save	[	239	]	;
				tuser_save	[	241	]	<=	tuser_save	[	240	]	;
				tuser_save	[	242	]	<=	tuser_save	[	241	]	;
				tuser_save	[	243	]	<=	tuser_save	[	242	]	;
				tuser_save	[	244	]	<=	tuser_save	[	243	]	;
				tuser_save	[	245	]	<=	tuser_save	[	244	]	;
				tuser_save	[	246	]	<=	tuser_save	[	245	]	;
				tuser_save	[	247	]	<=	tuser_save	[	246	]	;
				tuser_save	[	248	]	<=	tuser_save	[	247	]	;
				tuser_save	[	249	]	<=	tuser_save	[	248	]	;
				tuser_save	[	250	]	<=	tuser_save	[	249	]	;
				tuser_save	[	251	]	<=	tuser_save	[	250	]	;
				tuser_save	[	252	]	<=	tuser_save	[	251	]	;
				tuser_save	[	253	]	<=	tuser_save	[	252	]	;
				tuser_save	[	254	]	<=	tuser_save	[	253	]	;
				tuser_save	[	255	]	<=	tuser_save	[	254	]	;
					if(count_packet == 2'd2)
					begin
						count_packet <= 2'd0;
					end
					else
					begin
						count_packet	<= count_packet + 1'b1;
					end
					sum_tdata		<=	tdata_save[255];
					sum_tuser		<=	tuser_save[127];
					sum_tdata_valid		<=	1'b1;
					sum_tuser_valid		<=	1'b1;
				end
				else if(count_packet == 2'd1)
				begin
					tdata_save	[	0	]	<=	axififo_din;	//shift			
					tdata_save	[	1	]	<=	tdata_save	[	0	]	;
					tdata_save	[	2	]	<=	tdata_save	[	1	]	;
					tdata_save	[	3	]	<=	tdata_save	[	2	]	;
					tdata_save	[	4	]	<=	tdata_save	[	3	]	;
					tdata_save	[	5	]	<=	tdata_save	[	4	]	;
					tdata_save	[	6	]	<=	tdata_save	[	5	]	;
					tdata_save	[	7	]	<=	tdata_save	[	6	]	;
					tdata_save	[	8	]	<=	tdata_save	[	7	]	;
					tdata_save	[	9	]	<=	tdata_save	[	8	]	;
					tdata_save	[	10	]	<=	tdata_save	[	9	]	;
					tdata_save	[	11	]	<=	tdata_save	[	10	]	;
					tdata_save	[	12	]	<=	tdata_save	[	11	]	;
					tdata_save	[	13	]	<=	tdata_save	[	12	]	;
					tdata_save	[	14	]	<=	tdata_save	[	13	]	;
					tdata_save	[	15	]	<=	tdata_save	[	14	]	;
					tdata_save	[	16	]	<=	tdata_save	[	15	]	;
					tdata_save	[	17	]	<=	tdata_save	[	16	]	;
					tdata_save	[	18	]	<=	tdata_save	[	17	]	;
					tdata_save	[	19	]	<=	tdata_save	[	18	]	;
					tdata_save	[	20	]	<=	tdata_save	[	19	]	;
					tdata_save	[	21	]	<=	tdata_save	[	20	]	;
					tdata_save	[	22	]	<=	tdata_save	[	21	]	;
					tdata_save	[	23	]	<=	tdata_save	[	22	]	;
					tdata_save	[	24	]	<=	tdata_save	[	23	]	;
					tdata_save	[	25	]	<=	tdata_save	[	24	]	;
					tdata_save	[	26	]	<=	tdata_save	[	25	]	;
					tdata_save	[	27	]	<=	tdata_save	[	26	]	;
					tdata_save	[	28	]	<=	tdata_save	[	27	]	;
					tdata_save	[	29	]	<=	tdata_save	[	28	]	;
					tdata_save	[	30	]	<=	tdata_save	[	29	]	;
					tdata_save	[	31	]	<=	tdata_save	[	30	]	;
					tdata_save	[	32	]	<=	tdata_save	[	31	]	;
					tdata_save	[	33	]	<=	tdata_save	[	32	]	;
					tdata_save	[	34	]	<=	tdata_save	[	33	]	;
					tdata_save	[	35	]	<=	tdata_save	[	34	]	;
					tdata_save	[	36	]	<=	tdata_save	[	35	]	;
					tdata_save	[	37	]	<=	tdata_save	[	36	]	;
					tdata_save	[	38	]	<=	tdata_save	[	37	]	;
					tdata_save	[	39	]	<=	tdata_save	[	38	]	;
					tdata_save	[	40	]	<=	tdata_save	[	39	]	;
					tdata_save	[	41	]	<=	tdata_save	[	40	]	;
					tdata_save	[	42	]	<=	tdata_save	[	41	]	;
					tdata_save	[	43	]	<=	tdata_save	[	42	]	;
					tdata_save	[	44	]	<=	tdata_save	[	43	]	;
					tdata_save	[	45	]	<=	tdata_save	[	44	]	;
					tdata_save	[	46	]	<=	tdata_save	[	45	]	;
					tdata_save	[	47	]	<=	tdata_save	[	46	]	;
					tdata_save	[	48	]	<=	tdata_save	[	47	]	;
					tdata_save	[	49	]	<=	tdata_save	[	48	]	;
					tdata_save	[	50	]	<=	tdata_save	[	49	]	;
					tdata_save	[	51	]	<=	tdata_save	[	50	]	;
					tdata_save	[	52	]	<=	tdata_save	[	51	]	;
					tdata_save	[	53	]	<=	tdata_save	[	52	]	;
					tdata_save	[	54	]	<=	tdata_save	[	53	]	;
					tdata_save	[	55	]	<=	tdata_save	[	54	]	;
					tdata_save	[	56	]	<=	tdata_save	[	55	]	;
					tdata_save	[	57	]	<=	tdata_save	[	56	]	;
					tdata_save	[	58	]	<=	tdata_save	[	57	]	;
					tdata_save	[	59	]	<=	tdata_save	[	58	]	;
					tdata_save	[	60	]	<=	tdata_save	[	59	]	;
					tdata_save	[	61	]	<=	tdata_save	[	60	]	;
					tdata_save	[	62	]	<=	tdata_save	[	61	]	;
					tdata_save	[	63	]	<=	tdata_save	[	62	]	;
					tdata_save	[	64	]	<=	tdata_save	[	63	]	;
					tdata_save	[	65	]	<=	tdata_save	[	64	]	;
					tdata_save	[	66	]	<=	tdata_save	[	65	]	;
					tdata_save	[	67	]	<=	tdata_save	[	66	]	;
					tdata_save	[	68	]	<=	tdata_save	[	67	]	;
					tdata_save	[	69	]	<=	tdata_save	[	68	]	;
					tdata_save	[	70	]	<=	tdata_save	[	69	]	;
					tdata_save	[	71	]	<=	tdata_save	[	70	]	;
					tdata_save	[	72	]	<=	tdata_save	[	71	]	;
					tdata_save	[	73	]	<=	tdata_save	[	72	]	;
					tdata_save	[	74	]	<=	tdata_save	[	73	]	;
					tdata_save	[	75	]	<=	tdata_save	[	74	]	;
					tdata_save	[	76	]	<=	tdata_save	[	75	]	;
					tdata_save	[	77	]	<=	tdata_save	[	76	]	;
					tdata_save	[	78	]	<=	tdata_save	[	77	]	;
					tdata_save	[	79	]	<=	tdata_save	[	78	]	;
					tdata_save	[	80	]	<=	tdata_save	[	79	]	;
					tdata_save	[	81	]	<=	tdata_save	[	80	]	;
					tdata_save	[	82	]	<=	tdata_save	[	81	]	;
					tdata_save	[	83	]	<=	tdata_save	[	82	]	;
					tdata_save	[	84	]	<=	tdata_save	[	83	]	;
					tdata_save	[	85	]	<=	tdata_save	[	84	]	;
					tdata_save	[	86	]	<=	tdata_save	[	85	]	;
					tdata_save	[	87	]	<=	tdata_save	[	86	]	;
					tdata_save	[	88	]	<=	tdata_save	[	87	]	;
					tdata_save	[	89	]	<=	tdata_save	[	88	]	;
					tdata_save	[	90	]	<=	tdata_save	[	89	]	;
					tdata_save	[	91	]	<=	tdata_save	[	90	]	;
					tdata_save	[	92	]	<=	tdata_save	[	91	]	;
					tdata_save	[	93	]	<=	tdata_save	[	92	]	;
					tdata_save	[	94	]	<=	tdata_save	[	93	]	;
					tdata_save	[	95	]	<=	tdata_save	[	94	]	;
					tdata_save	[	96	]	<=	tdata_save	[	95	]	;
					tdata_save	[	97	]	<=	tdata_save	[	96	]	;
					tdata_save	[	98	]	<=	tdata_save	[	97	]	;
					tdata_save	[	99	]	<=	tdata_save	[	98	]	;
					tdata_save	[	100	]	<=	tdata_save	[	99	]	;
					tdata_save	[	101	]	<=	tdata_save	[	100	]	;
					tdata_save	[	102	]	<=	tdata_save	[	101	]	;
					tdata_save	[	103	]	<=	tdata_save	[	102	]	;
					tdata_save	[	104	]	<=	tdata_save	[	103	]	;
					tdata_save	[	105	]	<=	tdata_save	[	104	]	;
					tdata_save	[	106	]	<=	tdata_save	[	105	]	;
					tdata_save	[	107	]	<=	tdata_save	[	106	]	;
					tdata_save	[	108	]	<=	tdata_save	[	107	]	;
					tdata_save	[	109	]	<=	tdata_save	[	108	]	;
					tdata_save	[	110	]	<=	tdata_save	[	109	]	;
					tdata_save	[	111	]	<=	tdata_save	[	110	]	;
					tdata_save	[	112	]	<=	tdata_save	[	111	]	;
					tdata_save	[	113	]	<=	tdata_save	[	112	]	;
					tdata_save	[	114	]	<=	tdata_save	[	113	]	;
					tdata_save	[	115	]	<=	tdata_save	[	114	]	;
					tdata_save	[	116	]	<=	tdata_save	[	115	]	;
					tdata_save	[	117	]	<=	tdata_save	[	116	]	;
					tdata_save	[	118	]	<=	tdata_save	[	117	]	;
					tdata_save	[	119	]	<=	tdata_save	[	118	]	;
					tdata_save	[	120	]	<=	tdata_save	[	119	]	;
					tdata_save	[	121	]	<=	tdata_save	[	120	]	;
					tdata_save	[	122	]	<=	tdata_save	[	121	]	;
					tdata_save	[	123	]	<=	tdata_save	[	122	]	;
					tdata_save	[	124	]	<=	tdata_save	[	123	]	;
					tdata_save	[	125	]	<=	tdata_save	[	124	]	;
					tdata_save	[	126	]	<=	tdata_save	[	125	]	;
					tdata_save	[	127	]	<=	tdata_save	[	126	]	;
					tdata_save	[	128	]	<=	tdata_save	[	127	]	;
					tdata_save	[	129	]	<=	tdata_save	[	128	]	;
					tdata_save	[	130	]	<=	tdata_save	[	129	]	;
					tdata_save	[	131	]	<=	tdata_save	[	130	]	;
					tdata_save	[	132	]	<=	tdata_save	[	131	]	;
					tdata_save	[	133	]	<=	tdata_save	[	132	]	;
					tdata_save	[	134	]	<=	tdata_save	[	133	]	;
					tdata_save	[	135	]	<=	tdata_save	[	134	]	;
					tdata_save	[	136	]	<=	tdata_save	[	135	]	;
					tdata_save	[	137	]	<=	tdata_save	[	136	]	;
					tdata_save	[	138	]	<=	tdata_save	[	137	]	;
					tdata_save	[	139	]	<=	tdata_save	[	138	]	;
					tdata_save	[	140	]	<=	tdata_save	[	139	]	;
					tdata_save	[	141	]	<=	tdata_save	[	140	]	;
					tdata_save	[	142	]	<=	tdata_save	[	141	]	;
					tdata_save	[	143	]	<=	tdata_save	[	142	]	;
					tdata_save	[	144	]	<=	tdata_save	[	143	]	;
					tdata_save	[	145	]	<=	tdata_save	[	144	]	;
					tdata_save	[	146	]	<=	tdata_save	[	145	]	;
					tdata_save	[	147	]	<=	tdata_save	[	146	]	;
					tdata_save	[	148	]	<=	tdata_save	[	147	]	;
					tdata_save	[	149	]	<=	tdata_save	[	148	]	;
					tdata_save	[	150	]	<=	tdata_save	[	149	]	;
					tdata_save	[	151	]	<=	tdata_save	[	150	]	;
					tdata_save	[	152	]	<=	tdata_save	[	151	]	;
					tdata_save	[	153	]	<=	tdata_save	[	152	]	;
					tdata_save	[	154	]	<=	tdata_save	[	153	]	;
					tdata_save	[	155	]	<=	tdata_save	[	154	]	;
					tdata_save	[	156	]	<=	tdata_save	[	155	]	;
					tdata_save	[	157	]	<=	tdata_save	[	156	]	;
					tdata_save	[	158	]	<=	tdata_save	[	157	]	;
					tdata_save	[	159	]	<=	tdata_save	[	158	]	;
					tdata_save	[	160	]	<=	tdata_save	[	159	]	;
					tdata_save	[	161	]	<=	tdata_save	[	160	]	;
					tdata_save	[	162	]	<=	tdata_save	[	161	]	;
					tdata_save	[	163	]	<=	tdata_save	[	162	]	;
					tdata_save	[	164	]	<=	tdata_save	[	163	]	;
					tdata_save	[	165	]	<=	tdata_save	[	164	]	;
					tdata_save	[	166	]	<=	tdata_save	[	165	]	;
					tdata_save	[	167	]	<=	tdata_save	[	166	]	;
					tdata_save	[	168	]	<=	tdata_save	[	167	]	;
					tdata_save	[	169	]	<=	tdata_save	[	168	]	;
					tdata_save	[	170	]	<=	tdata_save	[	169	]	;
					tdata_save	[	171	]	<=	tdata_save	[	170	]	;
					tdata_save	[	172	]	<=	tdata_save	[	171	]	;
					tdata_save	[	173	]	<=	tdata_save	[	172	]	;
					tdata_save	[	174	]	<=	tdata_save	[	173	]	;
					tdata_save	[	175	]	<=	tdata_save	[	174	]	;
					tdata_save	[	176	]	<=	tdata_save	[	175	]	;
					tdata_save	[	177	]	<=	tdata_save	[	176	]	;
					tdata_save	[	178	]	<=	tdata_save	[	177	]	;
					tdata_save	[	179	]	<=	tdata_save	[	178	]	;
					tdata_save	[	180	]	<=	tdata_save	[	179	]	;
					tdata_save	[	181	]	<=	tdata_save	[	180	]	;
					tdata_save	[	182	]	<=	tdata_save	[	181	]	;
					tdata_save	[	183	]	<=	tdata_save	[	182	]	;
					tdata_save	[	184	]	<=	tdata_save	[	183	]	;
					tdata_save	[	185	]	<=	tdata_save	[	184	]	;
					tdata_save	[	186	]	<=	tdata_save	[	185	]	;
					tdata_save	[	187	]	<=	tdata_save	[	186	]	;
					tdata_save	[	188	]	<=	tdata_save	[	187	]	;
					tdata_save	[	189	]	<=	tdata_save	[	188	]	;
					tdata_save	[	190	]	<=	tdata_save	[	189	]	;
					tdata_save	[	191	]	<=	tdata_save	[	190	]	;
					tdata_save	[	192	]	<=	tdata_save	[	191	]	;
					tdata_save	[	193	]	<=	tdata_save	[	192	]	;
					tdata_save	[	194	]	<=	tdata_save	[	193	]	;
					tdata_save	[	195	]	<=	tdata_save	[	194	]	;
					tdata_save	[	196	]	<=	tdata_save	[	195	]	;
					tdata_save	[	197	]	<=	tdata_save	[	196	]	;
					tdata_save	[	198	]	<=	tdata_save	[	197	]	;
					tdata_save	[	199	]	<=	tdata_save	[	198	]	;
					tdata_save	[	200	]	<=	tdata_save	[	199	]	;
					tdata_save	[	201	]	<=	tdata_save	[	200	]	;
					tdata_save	[	202	]	<=	tdata_save	[	201	]	;
					tdata_save	[	203	]	<=	tdata_save	[	202	]	;
					tdata_save	[	204	]	<=	tdata_save	[	203	]	;
					tdata_save	[	205	]	<=	tdata_save	[	204	]	;
					tdata_save	[	206	]	<=	tdata_save	[	205	]	;
					tdata_save	[	207	]	<=	tdata_save	[	206	]	;
					tdata_save	[	208	]	<=	tdata_save	[	207	]	;
					tdata_save	[	209	]	<=	tdata_save	[	208	]	;
					tdata_save	[	210	]	<=	tdata_save	[	209	]	;
					tdata_save	[	211	]	<=	tdata_save	[	210	]	;
					tdata_save	[	212	]	<=	tdata_save	[	211	]	;
					tdata_save	[	213	]	<=	tdata_save	[	212	]	;
					tdata_save	[	214	]	<=	tdata_save	[	213	]	;
					tdata_save	[	215	]	<=	tdata_save	[	214	]	;
					tdata_save	[	216	]	<=	tdata_save	[	215	]	;
					tdata_save	[	217	]	<=	tdata_save	[	216	]	;
					tdata_save	[	218	]	<=	tdata_save	[	217	]	;
					tdata_save	[	219	]	<=	tdata_save	[	218	]	;
					tdata_save	[	220	]	<=	tdata_save	[	219	]	;
					tdata_save	[	221	]	<=	tdata_save	[	220	]	;
					tdata_save	[	222	]	<=	tdata_save	[	221	]	;
					tdata_save	[	223	]	<=	tdata_save	[	222	]	;
					tdata_save	[	224	]	<=	tdata_save	[	223	]	;
					tdata_save	[	225	]	<=	tdata_save	[	224	]	;
					tdata_save	[	226	]	<=	tdata_save	[	225	]	;
					tdata_save	[	227	]	<=	tdata_save	[	226	]	;
					tdata_save	[	228	]	<=	tdata_save	[	227	]	;
					tdata_save	[	229	]	<=	tdata_save	[	228	]	;
					tdata_save	[	230	]	<=	tdata_save	[	229	]	;
					tdata_save	[	231	]	<=	tdata_save	[	230	]	;
					tdata_save	[	232	]	<=	tdata_save	[	231	]	;
					tdata_save	[	233	]	<=	tdata_save	[	232	]	;
					tdata_save	[	234	]	<=	tdata_save	[	233	]	;
					tdata_save	[	235	]	<=	tdata_save	[	234	]	;
					tdata_save	[	236	]	<=	tdata_save	[	235	]	;
					tdata_save	[	237	]	<=	tdata_save	[	236	]	;
					tdata_save	[	238	]	<=	tdata_save	[	237	]	;
					tdata_save	[	239	]	<=	tdata_save	[	238	]	;
					tdata_save	[	240	]	<=	tdata_save	[	239	]	;
					tdata_save	[	241	]	<=	tdata_save	[	240	]	;
					tdata_save	[	242	]	<=	tdata_save	[	241	]	;
					tdata_save	[	243	]	<=	tdata_save	[	242	]	;
					tdata_save	[	244	]	<=	tdata_save	[	243	]	;
					tdata_save	[	245	]	<=	tdata_save	[	244	]	;
					tdata_save	[	246	]	<=	tdata_save	[	245	]	;
					tdata_save	[	247	]	<=	tdata_save	[	246	]	;
					tdata_save	[	248	]	<=	tdata_save	[	247	]	;
					tdata_save	[	249	]	<=	tdata_save	[	248	]	;
					tdata_save	[	250	]	<=	tdata_save	[	249	]	;
					tdata_save	[	251	]	<=	tdata_save	[	250	]	;
					tdata_save	[	252	]	<=	tdata_save	[	251	]	;
					tdata_save	[	253	]	<=	tdata_save	[	252	]	;
					tdata_save	[	254	]	<=	tdata_save	[	253	]	;
					tdata_save	[	255	]	<=	tdata_save	[	254	]	;
					tuser_save	[	0	]	<=	tuser;						
				tuser_save	[	1	]	<=	tuser_save	[	0	]	;
				tuser_save	[	2	]	<=	tuser_save	[	1	]	;
				tuser_save	[	3	]	<=	tuser_save	[	2	]	;
				tuser_save	[	4	]	<=	tuser_save	[	3	]	;
				tuser_save	[	5	]	<=	tuser_save	[	4	]	;
				tuser_save	[	6	]	<=	tuser_save	[	5	]	;
				tuser_save	[	7	]	<=	tuser_save	[	6	]	;
				tuser_save	[	8	]	<=	tuser_save	[	7	]	;
				tuser_save	[	9	]	<=	tuser_save	[	8	]	;
				tuser_save	[	10	]	<=	tuser_save	[	9	]	;
				tuser_save	[	11	]	<=	tuser_save	[	10	]	;
				tuser_save	[	12	]	<=	tuser_save	[	11	]	;
				tuser_save	[	13	]	<=	tuser_save	[	12	]	;
				tuser_save	[	14	]	<=	tuser_save	[	13	]	;
				tuser_save	[	15	]	<=	tuser_save	[	14	]	;
				tuser_save	[	16	]	<=	tuser_save	[	15	]	;
				tuser_save	[	17	]	<=	tuser_save	[	16	]	;
				tuser_save	[	18	]	<=	tuser_save	[	17	]	;
				tuser_save	[	19	]	<=	tuser_save	[	18	]	;
				tuser_save	[	20	]	<=	tuser_save	[	19	]	;
				tuser_save	[	21	]	<=	tuser_save	[	20	]	;
				tuser_save	[	22	]	<=	tuser_save	[	21	]	;
				tuser_save	[	23	]	<=	tuser_save	[	22	]	;
				tuser_save	[	24	]	<=	tuser_save	[	23	]	;
				tuser_save	[	25	]	<=	tuser_save	[	24	]	;
				tuser_save	[	26	]	<=	tuser_save	[	25	]	;
				tuser_save	[	27	]	<=	tuser_save	[	26	]	;
				tuser_save	[	28	]	<=	tuser_save	[	27	]	;
				tuser_save	[	29	]	<=	tuser_save	[	28	]	;
				tuser_save	[	30	]	<=	tuser_save	[	29	]	;
				tuser_save	[	31	]	<=	tuser_save	[	30	]	;
				tuser_save	[	32	]	<=	tuser_save	[	31	]	;
				tuser_save	[	33	]	<=	tuser_save	[	32	]	;
				tuser_save	[	34	]	<=	tuser_save	[	33	]	;
				tuser_save	[	35	]	<=	tuser_save	[	34	]	;
				tuser_save	[	36	]	<=	tuser_save	[	35	]	;
				tuser_save	[	37	]	<=	tuser_save	[	36	]	;
				tuser_save	[	38	]	<=	tuser_save	[	37	]	;
				tuser_save	[	39	]	<=	tuser_save	[	38	]	;
				tuser_save	[	40	]	<=	tuser_save	[	39	]	;
				tuser_save	[	41	]	<=	tuser_save	[	40	]	;
				tuser_save	[	42	]	<=	tuser_save	[	41	]	;
				tuser_save	[	43	]	<=	tuser_save	[	42	]	;
				tuser_save	[	44	]	<=	tuser_save	[	43	]	;
				tuser_save	[	45	]	<=	tuser_save	[	44	]	;
				tuser_save	[	46	]	<=	tuser_save	[	45	]	;
				tuser_save	[	47	]	<=	tuser_save	[	46	]	;
				tuser_save	[	48	]	<=	tuser_save	[	47	]	;
				tuser_save	[	49	]	<=	tuser_save	[	48	]	;
				tuser_save	[	50	]	<=	tuser_save	[	49	]	;
				tuser_save	[	51	]	<=	tuser_save	[	50	]	;
				tuser_save	[	52	]	<=	tuser_save	[	51	]	;
				tuser_save	[	53	]	<=	tuser_save	[	52	]	;
				tuser_save	[	54	]	<=	tuser_save	[	53	]	;
				tuser_save	[	55	]	<=	tuser_save	[	54	]	;
				tuser_save	[	56	]	<=	tuser_save	[	55	]	;
				tuser_save	[	57	]	<=	tuser_save	[	56	]	;
				tuser_save	[	58	]	<=	tuser_save	[	57	]	;
				tuser_save	[	59	]	<=	tuser_save	[	58	]	;
				tuser_save	[	60	]	<=	tuser_save	[	59	]	;
				tuser_save	[	61	]	<=	tuser_save	[	60	]	;
				tuser_save	[	62	]	<=	tuser_save	[	61	]	;
				tuser_save	[	63	]	<=	tuser_save	[	62	]	;
				tuser_save	[	64	]	<=	tuser_save	[	63	]	;
				tuser_save	[	65	]	<=	tuser_save	[	64	]	;
				tuser_save	[	66	]	<=	tuser_save	[	65	]	;
				tuser_save	[	67	]	<=	tuser_save	[	66	]	;
				tuser_save	[	68	]	<=	tuser_save	[	67	]	;
				tuser_save	[	69	]	<=	tuser_save	[	68	]	;
				tuser_save	[	70	]	<=	tuser_save	[	69	]	;
				tuser_save	[	71	]	<=	tuser_save	[	70	]	;
				tuser_save	[	72	]	<=	tuser_save	[	71	]	;
				tuser_save	[	73	]	<=	tuser_save	[	72	]	;
				tuser_save	[	74	]	<=	tuser_save	[	73	]	;
				tuser_save	[	75	]	<=	tuser_save	[	74	]	;
				tuser_save	[	76	]	<=	tuser_save	[	75	]	;
				tuser_save	[	77	]	<=	tuser_save	[	76	]	;
				tuser_save	[	78	]	<=	tuser_save	[	77	]	;
				tuser_save	[	79	]	<=	tuser_save	[	78	]	;
				tuser_save	[	80	]	<=	tuser_save	[	79	]	;
				tuser_save	[	81	]	<=	tuser_save	[	80	]	;
				tuser_save	[	82	]	<=	tuser_save	[	81	]	;
				tuser_save	[	83	]	<=	tuser_save	[	82	]	;
				tuser_save	[	84	]	<=	tuser_save	[	83	]	;
				tuser_save	[	85	]	<=	tuser_save	[	84	]	;
				tuser_save	[	86	]	<=	tuser_save	[	85	]	;
				tuser_save	[	87	]	<=	tuser_save	[	86	]	;
				tuser_save	[	88	]	<=	tuser_save	[	87	]	;
				tuser_save	[	89	]	<=	tuser_save	[	88	]	;
				tuser_save	[	90	]	<=	tuser_save	[	89	]	;
				tuser_save	[	91	]	<=	tuser_save	[	90	]	;
				tuser_save	[	92	]	<=	tuser_save	[	91	]	;
				tuser_save	[	93	]	<=	tuser_save	[	92	]	;
				tuser_save	[	94	]	<=	tuser_save	[	93	]	;
				tuser_save	[	95	]	<=	tuser_save	[	94	]	;
				tuser_save	[	96	]	<=	tuser_save	[	95	]	;
				tuser_save	[	97	]	<=	tuser_save	[	96	]	;
				tuser_save	[	98	]	<=	tuser_save	[	97	]	;
				tuser_save	[	99	]	<=	tuser_save	[	98	]	;
				tuser_save	[	100	]	<=	tuser_save	[	99	]	;
				tuser_save	[	101	]	<=	tuser_save	[	100	]	;
				tuser_save	[	102	]	<=	tuser_save	[	101	]	;
				tuser_save	[	103	]	<=	tuser_save	[	102	]	;
				tuser_save	[	104	]	<=	tuser_save	[	103	]	;
				tuser_save	[	105	]	<=	tuser_save	[	104	]	;
				tuser_save	[	106	]	<=	tuser_save	[	105	]	;
				tuser_save	[	107	]	<=	tuser_save	[	106	]	;
				tuser_save	[	108	]	<=	tuser_save	[	107	]	;
				tuser_save	[	109	]	<=	tuser_save	[	108	]	;
				tuser_save	[	110	]	<=	tuser_save	[	109	]	;
				tuser_save	[	111	]	<=	tuser_save	[	110	]	;
				tuser_save	[	112	]	<=	tuser_save	[	111	]	;
				tuser_save	[	113	]	<=	tuser_save	[	112	]	;
				tuser_save	[	114	]	<=	tuser_save	[	113	]	;
				tuser_save	[	115	]	<=	tuser_save	[	114	]	;
				tuser_save	[	116	]	<=	tuser_save	[	115	]	;
				tuser_save	[	117	]	<=	tuser_save	[	116	]	;
				tuser_save	[	118	]	<=	tuser_save	[	117	]	;
				tuser_save	[	119	]	<=	tuser_save	[	118	]	;
				tuser_save	[	120	]	<=	tuser_save	[	119	]	;
				tuser_save	[	121	]	<=	tuser_save	[	120	]	;
				tuser_save	[	122	]	<=	tuser_save	[	121	]	;
				tuser_save	[	123	]	<=	tuser_save	[	122	]	;
				tuser_save	[	124	]	<=	tuser_save	[	123	]	;
				tuser_save	[	125	]	<=	tuser_save	[	124	]	;
				tuser_save	[	126	]	<=	tuser_save	[	125	]	;
				tuser_save	[	127	]	<=	tuser_save	[	126	]	;
				tuser_save	[	128	]	<=	tuser_save	[	127	]	;
				tuser_save	[	129	]	<=	tuser_save	[	128	]	;
				tuser_save	[	130	]	<=	tuser_save	[	129	]	;
				tuser_save	[	131	]	<=	tuser_save	[	130	]	;
				tuser_save	[	132	]	<=	tuser_save	[	131	]	;
				tuser_save	[	133	]	<=	tuser_save	[	132	]	;
				tuser_save	[	134	]	<=	tuser_save	[	133	]	;
				tuser_save	[	135	]	<=	tuser_save	[	134	]	;
				tuser_save	[	136	]	<=	tuser_save	[	135	]	;
				tuser_save	[	137	]	<=	tuser_save	[	136	]	;
				tuser_save	[	138	]	<=	tuser_save	[	137	]	;
				tuser_save	[	139	]	<=	tuser_save	[	138	]	;
				tuser_save	[	140	]	<=	tuser_save	[	139	]	;
				tuser_save	[	141	]	<=	tuser_save	[	140	]	;
				tuser_save	[	142	]	<=	tuser_save	[	141	]	;
				tuser_save	[	143	]	<=	tuser_save	[	142	]	;
				tuser_save	[	144	]	<=	tuser_save	[	143	]	;
				tuser_save	[	145	]	<=	tuser_save	[	144	]	;
				tuser_save	[	146	]	<=	tuser_save	[	145	]	;
				tuser_save	[	147	]	<=	tuser_save	[	146	]	;
				tuser_save	[	148	]	<=	tuser_save	[	147	]	;
				tuser_save	[	149	]	<=	tuser_save	[	148	]	;
				tuser_save	[	150	]	<=	tuser_save	[	149	]	;
				tuser_save	[	151	]	<=	tuser_save	[	150	]	;
				tuser_save	[	152	]	<=	tuser_save	[	151	]	;
				tuser_save	[	153	]	<=	tuser_save	[	152	]	;
				tuser_save	[	154	]	<=	tuser_save	[	153	]	;
				tuser_save	[	155	]	<=	tuser_save	[	154	]	;
				tuser_save	[	156	]	<=	tuser_save	[	155	]	;
				tuser_save	[	157	]	<=	tuser_save	[	156	]	;
				tuser_save	[	158	]	<=	tuser_save	[	157	]	;
				tuser_save	[	159	]	<=	tuser_save	[	158	]	;
				tuser_save	[	160	]	<=	tuser_save	[	159	]	;
				tuser_save	[	161	]	<=	tuser_save	[	160	]	;
				tuser_save	[	162	]	<=	tuser_save	[	161	]	;
				tuser_save	[	163	]	<=	tuser_save	[	162	]	;
				tuser_save	[	164	]	<=	tuser_save	[	163	]	;
				tuser_save	[	165	]	<=	tuser_save	[	164	]	;
				tuser_save	[	166	]	<=	tuser_save	[	165	]	;
				tuser_save	[	167	]	<=	tuser_save	[	166	]	;
				tuser_save	[	168	]	<=	tuser_save	[	167	]	;
				tuser_save	[	169	]	<=	tuser_save	[	168	]	;
				tuser_save	[	170	]	<=	tuser_save	[	169	]	;
				tuser_save	[	171	]	<=	tuser_save	[	170	]	;
				tuser_save	[	172	]	<=	tuser_save	[	171	]	;
				tuser_save	[	173	]	<=	tuser_save	[	172	]	;
				tuser_save	[	174	]	<=	tuser_save	[	173	]	;
				tuser_save	[	175	]	<=	tuser_save	[	174	]	;
				tuser_save	[	176	]	<=	tuser_save	[	175	]	;
				tuser_save	[	177	]	<=	tuser_save	[	176	]	;
				tuser_save	[	178	]	<=	tuser_save	[	177	]	;
				tuser_save	[	179	]	<=	tuser_save	[	178	]	;
				tuser_save	[	180	]	<=	tuser_save	[	179	]	;
				tuser_save	[	181	]	<=	tuser_save	[	180	]	;
				tuser_save	[	182	]	<=	tuser_save	[	181	]	;
				tuser_save	[	183	]	<=	tuser_save	[	182	]	;
				tuser_save	[	184	]	<=	tuser_save	[	183	]	;
				tuser_save	[	185	]	<=	tuser_save	[	184	]	;
				tuser_save	[	186	]	<=	tuser_save	[	185	]	;
				tuser_save	[	187	]	<=	tuser_save	[	186	]	;
				tuser_save	[	188	]	<=	tuser_save	[	187	]	;
				tuser_save	[	189	]	<=	tuser_save	[	188	]	;
				tuser_save	[	190	]	<=	tuser_save	[	189	]	;
				tuser_save	[	191	]	<=	tuser_save	[	190	]	;
				tuser_save	[	192	]	<=	tuser_save	[	191	]	;
				tuser_save	[	193	]	<=	tuser_save	[	192	]	;
				tuser_save	[	194	]	<=	tuser_save	[	193	]	;
				tuser_save	[	195	]	<=	tuser_save	[	194	]	;
				tuser_save	[	196	]	<=	tuser_save	[	195	]	;
				tuser_save	[	197	]	<=	tuser_save	[	196	]	;
				tuser_save	[	198	]	<=	tuser_save	[	197	]	;
				tuser_save	[	199	]	<=	tuser_save	[	198	]	;
				tuser_save	[	200	]	<=	tuser_save	[	199	]	;
				tuser_save	[	201	]	<=	tuser_save	[	200	]	;
				tuser_save	[	202	]	<=	tuser_save	[	201	]	;
				tuser_save	[	203	]	<=	tuser_save	[	202	]	;
				tuser_save	[	204	]	<=	tuser_save	[	203	]	;
				tuser_save	[	205	]	<=	tuser_save	[	204	]	;
				tuser_save	[	206	]	<=	tuser_save	[	205	]	;
				tuser_save	[	207	]	<=	tuser_save	[	206	]	;
				tuser_save	[	208	]	<=	tuser_save	[	207	]	;
				tuser_save	[	209	]	<=	tuser_save	[	208	]	;
				tuser_save	[	210	]	<=	tuser_save	[	209	]	;
				tuser_save	[	211	]	<=	tuser_save	[	210	]	;
				tuser_save	[	212	]	<=	tuser_save	[	211	]	;
				tuser_save	[	213	]	<=	tuser_save	[	212	]	;
				tuser_save	[	214	]	<=	tuser_save	[	213	]	;
				tuser_save	[	215	]	<=	tuser_save	[	214	]	;
				tuser_save	[	216	]	<=	tuser_save	[	215	]	;
				tuser_save	[	217	]	<=	tuser_save	[	216	]	;
				tuser_save	[	218	]	<=	tuser_save	[	217	]	;
				tuser_save	[	219	]	<=	tuser_save	[	218	]	;
				tuser_save	[	220	]	<=	tuser_save	[	219	]	;
				tuser_save	[	221	]	<=	tuser_save	[	220	]	;
				tuser_save	[	222	]	<=	tuser_save	[	221	]	;
				tuser_save	[	223	]	<=	tuser_save	[	222	]	;
				tuser_save	[	224	]	<=	tuser_save	[	223	]	;
				tuser_save	[	225	]	<=	tuser_save	[	224	]	;
				tuser_save	[	226	]	<=	tuser_save	[	225	]	;
				tuser_save	[	227	]	<=	tuser_save	[	226	]	;
				tuser_save	[	228	]	<=	tuser_save	[	227	]	;
				tuser_save	[	229	]	<=	tuser_save	[	228	]	;
				tuser_save	[	230	]	<=	tuser_save	[	229	]	;
				tuser_save	[	231	]	<=	tuser_save	[	230	]	;
				tuser_save	[	232	]	<=	tuser_save	[	231	]	;
				tuser_save	[	233	]	<=	tuser_save	[	232	]	;
				tuser_save	[	234	]	<=	tuser_save	[	233	]	;
				tuser_save	[	235	]	<=	tuser_save	[	234	]	;
				tuser_save	[	236	]	<=	tuser_save	[	235	]	;
				tuser_save	[	237	]	<=	tuser_save	[	236	]	;
				tuser_save	[	238	]	<=	tuser_save	[	237	]	;
				tuser_save	[	239	]	<=	tuser_save	[	238	]	;
				tuser_save	[	240	]	<=	tuser_save	[	239	]	;
				tuser_save	[	241	]	<=	tuser_save	[	240	]	;
				tuser_save	[	242	]	<=	tuser_save	[	241	]	;
				tuser_save	[	243	]	<=	tuser_save	[	242	]	;
				tuser_save	[	244	]	<=	tuser_save	[	243	]	;
				tuser_save	[	245	]	<=	tuser_save	[	244	]	;
				tuser_save	[	246	]	<=	tuser_save	[	245	]	;
				tuser_save	[	247	]	<=	tuser_save	[	246	]	;
				tuser_save	[	248	]	<=	tuser_save	[	247	]	;
				tuser_save	[	249	]	<=	tuser_save	[	248	]	;
				tuser_save	[	250	]	<=	tuser_save	[	249	]	;
				tuser_save	[	251	]	<=	tuser_save	[	250	]	;
				tuser_save	[	252	]	<=	tuser_save	[	251	]	;
				tuser_save	[	253	]	<=	tuser_save	[	252	]	;
				tuser_save	[	254	]	<=	tuser_save	[	253	]	;
				tuser_save	[	255	]	<=	tuser_save	[	254	]	;
					if(count_packet == 2'd2)
					begin
						count_packet <= 2'd0;
					end
					else
					begin
						count_packet	<= count_packet + 1'b1;
					end
					sum_tdata		<=	tdata_save[255];
					sum_tuser		<=	tuser_save[127];
					sum_tdata_valid		<=	1'b1;
					sum_tuser_valid		<=	1'b1;
				end
				else
				begin				
					tdata_save	[	0	]	<=	201'd0;	//shift			
					tdata_save	[	1	]	<=	tdata_save	[	0	]	;
					tdata_save	[	2	]	<=	tdata_save	[	1	]	;
					tdata_save	[	3	]	<=	tdata_save	[	2	]	;
					tdata_save	[	4	]	<=	tdata_save	[	3	]	;
					tdata_save	[	5	]	<=	tdata_save	[	4	]	;
					tdata_save	[	6	]	<=	tdata_save	[	5	]	;
					tdata_save	[	7	]	<=	tdata_save	[	6	]	;
					tdata_save	[	8	]	<=	tdata_save	[	7	]	;
					tdata_save	[	9	]	<=	tdata_save	[	8	]	;
					tdata_save	[	10	]	<=	tdata_save	[	9	]	;
					tdata_save	[	11	]	<=	tdata_save	[	10	]	;
					tdata_save	[	12	]	<=	tdata_save	[	11	]	;
					tdata_save	[	13	]	<=	tdata_save	[	12	]	;
					tdata_save	[	14	]	<=	tdata_save	[	13	]	;
					tdata_save	[	15	]	<=	tdata_save	[	14	]	;
					tdata_save	[	16	]	<=	tdata_save	[	15	]	;
					tdata_save	[	17	]	<=	tdata_save	[	16	]	;
					tdata_save	[	18	]	<=	tdata_save	[	17	]	;
					tdata_save	[	19	]	<=	tdata_save	[	18	]	;
					tdata_save	[	20	]	<=	tdata_save	[	19	]	;
					tdata_save	[	21	]	<=	tdata_save	[	20	]	;
					tdata_save	[	22	]	<=	tdata_save	[	21	]	;
					tdata_save	[	23	]	<=	tdata_save	[	22	]	;
					tdata_save	[	24	]	<=	tdata_save	[	23	]	;
					tdata_save	[	25	]	<=	tdata_save	[	24	]	;
					tdata_save	[	26	]	<=	tdata_save	[	25	]	;
					tdata_save	[	27	]	<=	tdata_save	[	26	]	;
					tdata_save	[	28	]	<=	tdata_save	[	27	]	;
					tdata_save	[	29	]	<=	tdata_save	[	28	]	;
					tdata_save	[	30	]	<=	tdata_save	[	29	]	;
					tdata_save	[	31	]	<=	tdata_save	[	30	]	;
					tdata_save	[	32	]	<=	tdata_save	[	31	]	;
					tdata_save	[	33	]	<=	tdata_save	[	32	]	;
					tdata_save	[	34	]	<=	tdata_save	[	33	]	;
					tdata_save	[	35	]	<=	tdata_save	[	34	]	;
					tdata_save	[	36	]	<=	tdata_save	[	35	]	;
					tdata_save	[	37	]	<=	tdata_save	[	36	]	;
					tdata_save	[	38	]	<=	tdata_save	[	37	]	;
					tdata_save	[	39	]	<=	tdata_save	[	38	]	;
					tdata_save	[	40	]	<=	tdata_save	[	39	]	;
					tdata_save	[	41	]	<=	tdata_save	[	40	]	;
					tdata_save	[	42	]	<=	tdata_save	[	41	]	;
					tdata_save	[	43	]	<=	tdata_save	[	42	]	;
					tdata_save	[	44	]	<=	tdata_save	[	43	]	;
					tdata_save	[	45	]	<=	tdata_save	[	44	]	;
					tdata_save	[	46	]	<=	tdata_save	[	45	]	;
					tdata_save	[	47	]	<=	tdata_save	[	46	]	;
					tdata_save	[	48	]	<=	tdata_save	[	47	]	;
					tdata_save	[	49	]	<=	tdata_save	[	48	]	;
					tdata_save	[	50	]	<=	tdata_save	[	49	]	;
					tdata_save	[	51	]	<=	tdata_save	[	50	]	;
					tdata_save	[	52	]	<=	tdata_save	[	51	]	;
					tdata_save	[	53	]	<=	tdata_save	[	52	]	;
					tdata_save	[	54	]	<=	tdata_save	[	53	]	;
					tdata_save	[	55	]	<=	tdata_save	[	54	]	;
					tdata_save	[	56	]	<=	tdata_save	[	55	]	;
					tdata_save	[	57	]	<=	tdata_save	[	56	]	;
					tdata_save	[	58	]	<=	tdata_save	[	57	]	;
					tdata_save	[	59	]	<=	tdata_save	[	58	]	;
					tdata_save	[	60	]	<=	tdata_save	[	59	]	;
					tdata_save	[	61	]	<=	tdata_save	[	60	]	;
					tdata_save	[	62	]	<=	tdata_save	[	61	]	;
					tdata_save	[	63	]	<=	tdata_save	[	62	]	;
					tdata_save	[	64	]	<=	tdata_save	[	63	]	;
					tdata_save	[	65	]	<=	tdata_save	[	64	]	;
					tdata_save	[	66	]	<=	tdata_save	[	65	]	;
					tdata_save	[	67	]	<=	tdata_save	[	66	]	;
					tdata_save	[	68	]	<=	tdata_save	[	67	]	;
					tdata_save	[	69	]	<=	tdata_save	[	68	]	;
					tdata_save	[	70	]	<=	tdata_save	[	69	]	;
					tdata_save	[	71	]	<=	tdata_save	[	70	]	;
					tdata_save	[	72	]	<=	tdata_save	[	71	]	;
					tdata_save	[	73	]	<=	tdata_save	[	72	]	;
					tdata_save	[	74	]	<=	tdata_save	[	73	]	;
					tdata_save	[	75	]	<=	tdata_save	[	74	]	;
					tdata_save	[	76	]	<=	tdata_save	[	75	]	;
					tdata_save	[	77	]	<=	tdata_save	[	76	]	;
					tdata_save	[	78	]	<=	tdata_save	[	77	]	;
					tdata_save	[	79	]	<=	tdata_save	[	78	]	;
					tdata_save	[	80	]	<=	tdata_save	[	79	]	;
					tdata_save	[	81	]	<=	tdata_save	[	80	]	;
					tdata_save	[	82	]	<=	tdata_save	[	81	]	;
					tdata_save	[	83	]	<=	tdata_save	[	82	]	;
					tdata_save	[	84	]	<=	tdata_save	[	83	]	;
					tdata_save	[	85	]	<=	tdata_save	[	84	]	;
					tdata_save	[	86	]	<=	tdata_save	[	85	]	;
					tdata_save	[	87	]	<=	tdata_save	[	86	]	;
					tdata_save	[	88	]	<=	tdata_save	[	87	]	;
					tdata_save	[	89	]	<=	tdata_save	[	88	]	;
					tdata_save	[	90	]	<=	tdata_save	[	89	]	;
					tdata_save	[	91	]	<=	tdata_save	[	90	]	;
					tdata_save	[	92	]	<=	tdata_save	[	91	]	;
					tdata_save	[	93	]	<=	tdata_save	[	92	]	;
					tdata_save	[	94	]	<=	tdata_save	[	93	]	;
					tdata_save	[	95	]	<=	tdata_save	[	94	]	;
					tdata_save	[	96	]	<=	tdata_save	[	95	]	;
					tdata_save	[	97	]	<=	tdata_save	[	96	]	;
					tdata_save	[	98	]	<=	tdata_save	[	97	]	;
					tdata_save	[	99	]	<=	tdata_save	[	98	]	;
					tdata_save	[	100	]	<=	tdata_save	[	99	]	;
					tdata_save	[	101	]	<=	tdata_save	[	100	]	;
					tdata_save	[	102	]	<=	tdata_save	[	101	]	;
					tdata_save	[	103	]	<=	tdata_save	[	102	]	;
					tdata_save	[	104	]	<=	tdata_save	[	103	]	;
					tdata_save	[	105	]	<=	tdata_save	[	104	]	;
					tdata_save	[	106	]	<=	tdata_save	[	105	]	;
					tdata_save	[	107	]	<=	tdata_save	[	106	]	;
					tdata_save	[	108	]	<=	tdata_save	[	107	]	;
					tdata_save	[	109	]	<=	tdata_save	[	108	]	;
					tdata_save	[	110	]	<=	tdata_save	[	109	]	;
					tdata_save	[	111	]	<=	tdata_save	[	110	]	;
					tdata_save	[	112	]	<=	tdata_save	[	111	]	;
					tdata_save	[	113	]	<=	tdata_save	[	112	]	;
					tdata_save	[	114	]	<=	tdata_save	[	113	]	;
					tdata_save	[	115	]	<=	tdata_save	[	114	]	;
					tdata_save	[	116	]	<=	tdata_save	[	115	]	;
					tdata_save	[	117	]	<=	tdata_save	[	116	]	;
					tdata_save	[	118	]	<=	tdata_save	[	117	]	;
					tdata_save	[	119	]	<=	tdata_save	[	118	]	;
					tdata_save	[	120	]	<=	tdata_save	[	119	]	;
					tdata_save	[	121	]	<=	tdata_save	[	120	]	;
					tdata_save	[	122	]	<=	tdata_save	[	121	]	;
					tdata_save	[	123	]	<=	tdata_save	[	122	]	;
					tdata_save	[	124	]	<=	tdata_save	[	123	]	;
					tdata_save	[	125	]	<=	tdata_save	[	124	]	;
					tdata_save	[	126	]	<=	tdata_save	[	125	]	;
					tdata_save	[	127	]	<=	tdata_save	[	126	]	;
					tdata_save	[	128	]	<=	tdata_save	[	127	]	;
					tdata_save	[	129	]	<=	tdata_save	[	128	]	;
					tdata_save	[	130	]	<=	tdata_save	[	129	]	;
					tdata_save	[	131	]	<=	tdata_save	[	130	]	;
					tdata_save	[	132	]	<=	tdata_save	[	131	]	;
					tdata_save	[	133	]	<=	tdata_save	[	132	]	;
					tdata_save	[	134	]	<=	tdata_save	[	133	]	;
					tdata_save	[	135	]	<=	tdata_save	[	134	]	;
					tdata_save	[	136	]	<=	tdata_save	[	135	]	;
					tdata_save	[	137	]	<=	tdata_save	[	136	]	;
					tdata_save	[	138	]	<=	tdata_save	[	137	]	;
					tdata_save	[	139	]	<=	tdata_save	[	138	]	;
					tdata_save	[	140	]	<=	tdata_save	[	139	]	;
					tdata_save	[	141	]	<=	tdata_save	[	140	]	;
					tdata_save	[	142	]	<=	tdata_save	[	141	]	;
					tdata_save	[	143	]	<=	tdata_save	[	142	]	;
					tdata_save	[	144	]	<=	tdata_save	[	143	]	;
					tdata_save	[	145	]	<=	tdata_save	[	144	]	;
					tdata_save	[	146	]	<=	tdata_save	[	145	]	;
					tdata_save	[	147	]	<=	tdata_save	[	146	]	;
					tdata_save	[	148	]	<=	tdata_save	[	147	]	;
					tdata_save	[	149	]	<=	tdata_save	[	148	]	;
					tdata_save	[	150	]	<=	tdata_save	[	149	]	;
					tdata_save	[	151	]	<=	tdata_save	[	150	]	;
					tdata_save	[	152	]	<=	tdata_save	[	151	]	;
					tdata_save	[	153	]	<=	tdata_save	[	152	]	;
					tdata_save	[	154	]	<=	tdata_save	[	153	]	;
					tdata_save	[	155	]	<=	tdata_save	[	154	]	;
					tdata_save	[	156	]	<=	tdata_save	[	155	]	;
					tdata_save	[	157	]	<=	tdata_save	[	156	]	;
					tdata_save	[	158	]	<=	tdata_save	[	157	]	;
					tdata_save	[	159	]	<=	tdata_save	[	158	]	;
					tdata_save	[	160	]	<=	tdata_save	[	159	]	;
					tdata_save	[	161	]	<=	tdata_save	[	160	]	;
					tdata_save	[	162	]	<=	tdata_save	[	161	]	;
					tdata_save	[	163	]	<=	tdata_save	[	162	]	;
					tdata_save	[	164	]	<=	tdata_save	[	163	]	;
					tdata_save	[	165	]	<=	tdata_save	[	164	]	;
					tdata_save	[	166	]	<=	tdata_save	[	165	]	;
					tdata_save	[	167	]	<=	tdata_save	[	166	]	;
					tdata_save	[	168	]	<=	tdata_save	[	167	]	;
					tdata_save	[	169	]	<=	tdata_save	[	168	]	;
					tdata_save	[	170	]	<=	tdata_save	[	169	]	;
					tdata_save	[	171	]	<=	tdata_save	[	170	]	;
					tdata_save	[	172	]	<=	tdata_save	[	171	]	;
					tdata_save	[	173	]	<=	tdata_save	[	172	]	;
					tdata_save	[	174	]	<=	tdata_save	[	173	]	;
					tdata_save	[	175	]	<=	tdata_save	[	174	]	;
					tdata_save	[	176	]	<=	tdata_save	[	175	]	;
					tdata_save	[	177	]	<=	tdata_save	[	176	]	;
					tdata_save	[	178	]	<=	tdata_save	[	177	]	;
					tdata_save	[	179	]	<=	tdata_save	[	178	]	;
					tdata_save	[	180	]	<=	tdata_save	[	179	]	;
					tdata_save	[	181	]	<=	tdata_save	[	180	]	;
					tdata_save	[	182	]	<=	tdata_save	[	181	]	;
					tdata_save	[	183	]	<=	tdata_save	[	182	]	;
					tdata_save	[	184	]	<=	tdata_save	[	183	]	;
					tdata_save	[	185	]	<=	tdata_save	[	184	]	;
					tdata_save	[	186	]	<=	tdata_save	[	185	]	;
					tdata_save	[	187	]	<=	tdata_save	[	186	]	;
					tdata_save	[	188	]	<=	tdata_save	[	187	]	;
					tdata_save	[	189	]	<=	tdata_save	[	188	]	;
					tdata_save	[	190	]	<=	tdata_save	[	189	]	;
					tdata_save	[	191	]	<=	tdata_save	[	190	]	;
					tdata_save	[	192	]	<=	tdata_save	[	191	]	;
					tdata_save	[	193	]	<=	tdata_save	[	192	]	;
					tdata_save	[	194	]	<=	tdata_save	[	193	]	;
					tdata_save	[	195	]	<=	tdata_save	[	194	]	;
					tdata_save	[	196	]	<=	tdata_save	[	195	]	;
					tdata_save	[	197	]	<=	tdata_save	[	196	]	;
					tdata_save	[	198	]	<=	tdata_save	[	197	]	;
					tdata_save	[	199	]	<=	tdata_save	[	198	]	;
					tdata_save	[	200	]	<=	tdata_save	[	199	]	;
					tdata_save	[	201	]	<=	tdata_save	[	200	]	;
					tdata_save	[	202	]	<=	tdata_save	[	201	]	;
					tdata_save	[	203	]	<=	tdata_save	[	202	]	;
					tdata_save	[	204	]	<=	tdata_save	[	203	]	;
					tdata_save	[	205	]	<=	tdata_save	[	204	]	;
					tdata_save	[	206	]	<=	tdata_save	[	205	]	;
					tdata_save	[	207	]	<=	tdata_save	[	206	]	;
					tdata_save	[	208	]	<=	tdata_save	[	207	]	;
					tdata_save	[	209	]	<=	tdata_save	[	208	]	;
					tdata_save	[	210	]	<=	tdata_save	[	209	]	;
					tdata_save	[	211	]	<=	tdata_save	[	210	]	;
					tdata_save	[	212	]	<=	tdata_save	[	211	]	;
					tdata_save	[	213	]	<=	tdata_save	[	212	]	;
					tdata_save	[	214	]	<=	tdata_save	[	213	]	;
					tdata_save	[	215	]	<=	tdata_save	[	214	]	;
					tdata_save	[	216	]	<=	tdata_save	[	215	]	;
					tdata_save	[	217	]	<=	tdata_save	[	216	]	;
					tdata_save	[	218	]	<=	tdata_save	[	217	]	;
					tdata_save	[	219	]	<=	tdata_save	[	218	]	;
					tdata_save	[	220	]	<=	tdata_save	[	219	]	;
					tdata_save	[	221	]	<=	tdata_save	[	220	]	;
					tdata_save	[	222	]	<=	tdata_save	[	221	]	;
					tdata_save	[	223	]	<=	tdata_save	[	222	]	;
					tdata_save	[	224	]	<=	tdata_save	[	223	]	;
					tdata_save	[	225	]	<=	tdata_save	[	224	]	;
					tdata_save	[	226	]	<=	tdata_save	[	225	]	;
					tdata_save	[	227	]	<=	tdata_save	[	226	]	;
					tdata_save	[	228	]	<=	tdata_save	[	227	]	;
					tdata_save	[	229	]	<=	tdata_save	[	228	]	;
					tdata_save	[	230	]	<=	tdata_save	[	229	]	;
					tdata_save	[	231	]	<=	tdata_save	[	230	]	;
					tdata_save	[	232	]	<=	tdata_save	[	231	]	;
					tdata_save	[	233	]	<=	tdata_save	[	232	]	;
					tdata_save	[	234	]	<=	tdata_save	[	233	]	;
					tdata_save	[	235	]	<=	tdata_save	[	234	]	;
					tdata_save	[	236	]	<=	tdata_save	[	235	]	;
					tdata_save	[	237	]	<=	tdata_save	[	236	]	;
					tdata_save	[	238	]	<=	tdata_save	[	237	]	;
					tdata_save	[	239	]	<=	tdata_save	[	238	]	;
					tdata_save	[	240	]	<=	tdata_save	[	239	]	;
					tdata_save	[	241	]	<=	tdata_save	[	240	]	;
					tdata_save	[	242	]	<=	tdata_save	[	241	]	;
					tdata_save	[	243	]	<=	tdata_save	[	242	]	;
					tdata_save	[	244	]	<=	tdata_save	[	243	]	;
					tdata_save	[	245	]	<=	tdata_save	[	244	]	;
					tdata_save	[	246	]	<=	tdata_save	[	245	]	;
					tdata_save	[	247	]	<=	tdata_save	[	246	]	;
					tdata_save	[	248	]	<=	tdata_save	[	247	]	;
					tdata_save	[	249	]	<=	tdata_save	[	248	]	;
					tdata_save	[	250	]	<=	tdata_save	[	249	]	;
					tdata_save	[	251	]	<=	tdata_save	[	250	]	;
					tdata_save	[	252	]	<=	tdata_save	[	251	]	;
					tdata_save	[	253	]	<=	tdata_save	[	252	]	;
					tdata_save	[	254	]	<=	tdata_save	[	253	]	;
					tdata_save	[	255	]	<=	tdata_save	[	254	]	;
					tuser_save	[	0	]	<=	128'd0;										
				tuser_save	[	1	]	<=	tuser_save	[	0	]	;
				tuser_save	[	2	]	<=	tuser_save	[	1	]	;
				tuser_save	[	3	]	<=	tuser_save	[	2	]	;
				tuser_save	[	4	]	<=	tuser_save	[	3	]	;
				tuser_save	[	5	]	<=	tuser_save	[	4	]	;
				tuser_save	[	6	]	<=	tuser_save	[	5	]	;
				tuser_save	[	7	]	<=	tuser_save	[	6	]	;
				tuser_save	[	8	]	<=	tuser_save	[	7	]	;
				tuser_save	[	9	]	<=	tuser_save	[	8	]	;
				tuser_save	[	10	]	<=	tuser_save	[	9	]	;
				tuser_save	[	11	]	<=	tuser_save	[	10	]	;
				tuser_save	[	12	]	<=	tuser_save	[	11	]	;
				tuser_save	[	13	]	<=	tuser_save	[	12	]	;
				tuser_save	[	14	]	<=	tuser_save	[	13	]	;
				tuser_save	[	15	]	<=	tuser_save	[	14	]	;
				tuser_save	[	16	]	<=	tuser_save	[	15	]	;
				tuser_save	[	17	]	<=	tuser_save	[	16	]	;
				tuser_save	[	18	]	<=	tuser_save	[	17	]	;
				tuser_save	[	19	]	<=	tuser_save	[	18	]	;
				tuser_save	[	20	]	<=	tuser_save	[	19	]	;
				tuser_save	[	21	]	<=	tuser_save	[	20	]	;
				tuser_save	[	22	]	<=	tuser_save	[	21	]	;
				tuser_save	[	23	]	<=	tuser_save	[	22	]	;
				tuser_save	[	24	]	<=	tuser_save	[	23	]	;
				tuser_save	[	25	]	<=	tuser_save	[	24	]	;
				tuser_save	[	26	]	<=	tuser_save	[	25	]	;
				tuser_save	[	27	]	<=	tuser_save	[	26	]	;
				tuser_save	[	28	]	<=	tuser_save	[	27	]	;
				tuser_save	[	29	]	<=	tuser_save	[	28	]	;
				tuser_save	[	30	]	<=	tuser_save	[	29	]	;
				tuser_save	[	31	]	<=	tuser_save	[	30	]	;
				tuser_save	[	32	]	<=	tuser_save	[	31	]	;
				tuser_save	[	33	]	<=	tuser_save	[	32	]	;
				tuser_save	[	34	]	<=	tuser_save	[	33	]	;
				tuser_save	[	35	]	<=	tuser_save	[	34	]	;
				tuser_save	[	36	]	<=	tuser_save	[	35	]	;
				tuser_save	[	37	]	<=	tuser_save	[	36	]	;
				tuser_save	[	38	]	<=	tuser_save	[	37	]	;
				tuser_save	[	39	]	<=	tuser_save	[	38	]	;
				tuser_save	[	40	]	<=	tuser_save	[	39	]	;
				tuser_save	[	41	]	<=	tuser_save	[	40	]	;
				tuser_save	[	42	]	<=	tuser_save	[	41	]	;
				tuser_save	[	43	]	<=	tuser_save	[	42	]	;
				tuser_save	[	44	]	<=	tuser_save	[	43	]	;
				tuser_save	[	45	]	<=	tuser_save	[	44	]	;
				tuser_save	[	46	]	<=	tuser_save	[	45	]	;
				tuser_save	[	47	]	<=	tuser_save	[	46	]	;
				tuser_save	[	48	]	<=	tuser_save	[	47	]	;
				tuser_save	[	49	]	<=	tuser_save	[	48	]	;
				tuser_save	[	50	]	<=	tuser_save	[	49	]	;
				tuser_save	[	51	]	<=	tuser_save	[	50	]	;
				tuser_save	[	52	]	<=	tuser_save	[	51	]	;
				tuser_save	[	53	]	<=	tuser_save	[	52	]	;
				tuser_save	[	54	]	<=	tuser_save	[	53	]	;
				tuser_save	[	55	]	<=	tuser_save	[	54	]	;
				tuser_save	[	56	]	<=	tuser_save	[	55	]	;
				tuser_save	[	57	]	<=	tuser_save	[	56	]	;
				tuser_save	[	58	]	<=	tuser_save	[	57	]	;
				tuser_save	[	59	]	<=	tuser_save	[	58	]	;
				tuser_save	[	60	]	<=	tuser_save	[	59	]	;
				tuser_save	[	61	]	<=	tuser_save	[	60	]	;
				tuser_save	[	62	]	<=	tuser_save	[	61	]	;
				tuser_save	[	63	]	<=	tuser_save	[	62	]	;
				tuser_save	[	64	]	<=	tuser_save	[	63	]	;
				tuser_save	[	65	]	<=	tuser_save	[	64	]	;
				tuser_save	[	66	]	<=	tuser_save	[	65	]	;
				tuser_save	[	67	]	<=	tuser_save	[	66	]	;
				tuser_save	[	68	]	<=	tuser_save	[	67	]	;
				tuser_save	[	69	]	<=	tuser_save	[	68	]	;
				tuser_save	[	70	]	<=	tuser_save	[	69	]	;
				tuser_save	[	71	]	<=	tuser_save	[	70	]	;
				tuser_save	[	72	]	<=	tuser_save	[	71	]	;
				tuser_save	[	73	]	<=	tuser_save	[	72	]	;
				tuser_save	[	74	]	<=	tuser_save	[	73	]	;
				tuser_save	[	75	]	<=	tuser_save	[	74	]	;
				tuser_save	[	76	]	<=	tuser_save	[	75	]	;
				tuser_save	[	77	]	<=	tuser_save	[	76	]	;
				tuser_save	[	78	]	<=	tuser_save	[	77	]	;
				tuser_save	[	79	]	<=	tuser_save	[	78	]	;
				tuser_save	[	80	]	<=	tuser_save	[	79	]	;
				tuser_save	[	81	]	<=	tuser_save	[	80	]	;
				tuser_save	[	82	]	<=	tuser_save	[	81	]	;
				tuser_save	[	83	]	<=	tuser_save	[	82	]	;
				tuser_save	[	84	]	<=	tuser_save	[	83	]	;
				tuser_save	[	85	]	<=	tuser_save	[	84	]	;
				tuser_save	[	86	]	<=	tuser_save	[	85	]	;
				tuser_save	[	87	]	<=	tuser_save	[	86	]	;
				tuser_save	[	88	]	<=	tuser_save	[	87	]	;
				tuser_save	[	89	]	<=	tuser_save	[	88	]	;
				tuser_save	[	90	]	<=	tuser_save	[	89	]	;
				tuser_save	[	91	]	<=	tuser_save	[	90	]	;
				tuser_save	[	92	]	<=	tuser_save	[	91	]	;
				tuser_save	[	93	]	<=	tuser_save	[	92	]	;
				tuser_save	[	94	]	<=	tuser_save	[	93	]	;
				tuser_save	[	95	]	<=	tuser_save	[	94	]	;
				tuser_save	[	96	]	<=	tuser_save	[	95	]	;
				tuser_save	[	97	]	<=	tuser_save	[	96	]	;
				tuser_save	[	98	]	<=	tuser_save	[	97	]	;
				tuser_save	[	99	]	<=	tuser_save	[	98	]	;
				tuser_save	[	100	]	<=	tuser_save	[	99	]	;
				tuser_save	[	101	]	<=	tuser_save	[	100	]	;
				tuser_save	[	102	]	<=	tuser_save	[	101	]	;
				tuser_save	[	103	]	<=	tuser_save	[	102	]	;
				tuser_save	[	104	]	<=	tuser_save	[	103	]	;
				tuser_save	[	105	]	<=	tuser_save	[	104	]	;
				tuser_save	[	106	]	<=	tuser_save	[	105	]	;
				tuser_save	[	107	]	<=	tuser_save	[	106	]	;
				tuser_save	[	108	]	<=	tuser_save	[	107	]	;
				tuser_save	[	109	]	<=	tuser_save	[	108	]	;
				tuser_save	[	110	]	<=	tuser_save	[	109	]	;
				tuser_save	[	111	]	<=	tuser_save	[	110	]	;
				tuser_save	[	112	]	<=	tuser_save	[	111	]	;
				tuser_save	[	113	]	<=	tuser_save	[	112	]	;
				tuser_save	[	114	]	<=	tuser_save	[	113	]	;
				tuser_save	[	115	]	<=	tuser_save	[	114	]	;
				tuser_save	[	116	]	<=	tuser_save	[	115	]	;
				tuser_save	[	117	]	<=	tuser_save	[	116	]	;
				tuser_save	[	118	]	<=	tuser_save	[	117	]	;
				tuser_save	[	119	]	<=	tuser_save	[	118	]	;
				tuser_save	[	120	]	<=	tuser_save	[	119	]	;
				tuser_save	[	121	]	<=	tuser_save	[	120	]	;
				tuser_save	[	122	]	<=	tuser_save	[	121	]	;
				tuser_save	[	123	]	<=	tuser_save	[	122	]	;
				tuser_save	[	124	]	<=	tuser_save	[	123	]	;
				tuser_save	[	125	]	<=	tuser_save	[	124	]	;
				tuser_save	[	126	]	<=	tuser_save	[	125	]	;
				tuser_save	[	127	]	<=	tuser_save	[	126	]	;
				tuser_save	[	128	]	<=	tuser_save	[	127	]	;
				tuser_save	[	129	]	<=	tuser_save	[	128	]	;
				tuser_save	[	130	]	<=	tuser_save	[	129	]	;
				tuser_save	[	131	]	<=	tuser_save	[	130	]	;
				tuser_save	[	132	]	<=	tuser_save	[	131	]	;
				tuser_save	[	133	]	<=	tuser_save	[	132	]	;
				tuser_save	[	134	]	<=	tuser_save	[	133	]	;
				tuser_save	[	135	]	<=	tuser_save	[	134	]	;
				tuser_save	[	136	]	<=	tuser_save	[	135	]	;
				tuser_save	[	137	]	<=	tuser_save	[	136	]	;
				tuser_save	[	138	]	<=	tuser_save	[	137	]	;
				tuser_save	[	139	]	<=	tuser_save	[	138	]	;
				tuser_save	[	140	]	<=	tuser_save	[	139	]	;
				tuser_save	[	141	]	<=	tuser_save	[	140	]	;
				tuser_save	[	142	]	<=	tuser_save	[	141	]	;
				tuser_save	[	143	]	<=	tuser_save	[	142	]	;
				tuser_save	[	144	]	<=	tuser_save	[	143	]	;
				tuser_save	[	145	]	<=	tuser_save	[	144	]	;
				tuser_save	[	146	]	<=	tuser_save	[	145	]	;
				tuser_save	[	147	]	<=	tuser_save	[	146	]	;
				tuser_save	[	148	]	<=	tuser_save	[	147	]	;
				tuser_save	[	149	]	<=	tuser_save	[	148	]	;
				tuser_save	[	150	]	<=	tuser_save	[	149	]	;
				tuser_save	[	151	]	<=	tuser_save	[	150	]	;
				tuser_save	[	152	]	<=	tuser_save	[	151	]	;
				tuser_save	[	153	]	<=	tuser_save	[	152	]	;
				tuser_save	[	154	]	<=	tuser_save	[	153	]	;
				tuser_save	[	155	]	<=	tuser_save	[	154	]	;
				tuser_save	[	156	]	<=	tuser_save	[	155	]	;
				tuser_save	[	157	]	<=	tuser_save	[	156	]	;
				tuser_save	[	158	]	<=	tuser_save	[	157	]	;
				tuser_save	[	159	]	<=	tuser_save	[	158	]	;
				tuser_save	[	160	]	<=	tuser_save	[	159	]	;
				tuser_save	[	161	]	<=	tuser_save	[	160	]	;
				tuser_save	[	162	]	<=	tuser_save	[	161	]	;
				tuser_save	[	163	]	<=	tuser_save	[	162	]	;
				tuser_save	[	164	]	<=	tuser_save	[	163	]	;
				tuser_save	[	165	]	<=	tuser_save	[	164	]	;
				tuser_save	[	166	]	<=	tuser_save	[	165	]	;
				tuser_save	[	167	]	<=	tuser_save	[	166	]	;
				tuser_save	[	168	]	<=	tuser_save	[	167	]	;
				tuser_save	[	169	]	<=	tuser_save	[	168	]	;
				tuser_save	[	170	]	<=	tuser_save	[	169	]	;
				tuser_save	[	171	]	<=	tuser_save	[	170	]	;
				tuser_save	[	172	]	<=	tuser_save	[	171	]	;
				tuser_save	[	173	]	<=	tuser_save	[	172	]	;
				tuser_save	[	174	]	<=	tuser_save	[	173	]	;
				tuser_save	[	175	]	<=	tuser_save	[	174	]	;
				tuser_save	[	176	]	<=	tuser_save	[	175	]	;
				tuser_save	[	177	]	<=	tuser_save	[	176	]	;
				tuser_save	[	178	]	<=	tuser_save	[	177	]	;
				tuser_save	[	179	]	<=	tuser_save	[	178	]	;
				tuser_save	[	180	]	<=	tuser_save	[	179	]	;
				tuser_save	[	181	]	<=	tuser_save	[	180	]	;
				tuser_save	[	182	]	<=	tuser_save	[	181	]	;
				tuser_save	[	183	]	<=	tuser_save	[	182	]	;
				tuser_save	[	184	]	<=	tuser_save	[	183	]	;
				tuser_save	[	185	]	<=	tuser_save	[	184	]	;
				tuser_save	[	186	]	<=	tuser_save	[	185	]	;
				tuser_save	[	187	]	<=	tuser_save	[	186	]	;
				tuser_save	[	188	]	<=	tuser_save	[	187	]	;
				tuser_save	[	189	]	<=	tuser_save	[	188	]	;
				tuser_save	[	190	]	<=	tuser_save	[	189	]	;
				tuser_save	[	191	]	<=	tuser_save	[	190	]	;
				tuser_save	[	192	]	<=	tuser_save	[	191	]	;
				tuser_save	[	193	]	<=	tuser_save	[	192	]	;
				tuser_save	[	194	]	<=	tuser_save	[	193	]	;
				tuser_save	[	195	]	<=	tuser_save	[	194	]	;
				tuser_save	[	196	]	<=	tuser_save	[	195	]	;
				tuser_save	[	197	]	<=	tuser_save	[	196	]	;
				tuser_save	[	198	]	<=	tuser_save	[	197	]	;
				tuser_save	[	199	]	<=	tuser_save	[	198	]	;
				tuser_save	[	200	]	<=	tuser_save	[	199	]	;
				tuser_save	[	201	]	<=	tuser_save	[	200	]	;
				tuser_save	[	202	]	<=	tuser_save	[	201	]	;
				tuser_save	[	203	]	<=	tuser_save	[	202	]	;
				tuser_save	[	204	]	<=	tuser_save	[	203	]	;
				tuser_save	[	205	]	<=	tuser_save	[	204	]	;
				tuser_save	[	206	]	<=	tuser_save	[	205	]	;
				tuser_save	[	207	]	<=	tuser_save	[	206	]	;
				tuser_save	[	208	]	<=	tuser_save	[	207	]	;
				tuser_save	[	209	]	<=	tuser_save	[	208	]	;
				tuser_save	[	210	]	<=	tuser_save	[	209	]	;
				tuser_save	[	211	]	<=	tuser_save	[	210	]	;
				tuser_save	[	212	]	<=	tuser_save	[	211	]	;
				tuser_save	[	213	]	<=	tuser_save	[	212	]	;
				tuser_save	[	214	]	<=	tuser_save	[	213	]	;
				tuser_save	[	215	]	<=	tuser_save	[	214	]	;
				tuser_save	[	216	]	<=	tuser_save	[	215	]	;
				tuser_save	[	217	]	<=	tuser_save	[	216	]	;
				tuser_save	[	218	]	<=	tuser_save	[	217	]	;
				tuser_save	[	219	]	<=	tuser_save	[	218	]	;
				tuser_save	[	220	]	<=	tuser_save	[	219	]	;
				tuser_save	[	221	]	<=	tuser_save	[	220	]	;
				tuser_save	[	222	]	<=	tuser_save	[	221	]	;
				tuser_save	[	223	]	<=	tuser_save	[	222	]	;
				tuser_save	[	224	]	<=	tuser_save	[	223	]	;
				tuser_save	[	225	]	<=	tuser_save	[	224	]	;
				tuser_save	[	226	]	<=	tuser_save	[	225	]	;
				tuser_save	[	227	]	<=	tuser_save	[	226	]	;
				tuser_save	[	228	]	<=	tuser_save	[	227	]	;
				tuser_save	[	229	]	<=	tuser_save	[	228	]	;
				tuser_save	[	230	]	<=	tuser_save	[	229	]	;
				tuser_save	[	231	]	<=	tuser_save	[	230	]	;
				tuser_save	[	232	]	<=	tuser_save	[	231	]	;
				tuser_save	[	233	]	<=	tuser_save	[	232	]	;
				tuser_save	[	234	]	<=	tuser_save	[	233	]	;
				tuser_save	[	235	]	<=	tuser_save	[	234	]	;
				tuser_save	[	236	]	<=	tuser_save	[	235	]	;
				tuser_save	[	237	]	<=	tuser_save	[	236	]	;
				tuser_save	[	238	]	<=	tuser_save	[	237	]	;
				tuser_save	[	239	]	<=	tuser_save	[	238	]	;
				tuser_save	[	240	]	<=	tuser_save	[	239	]	;
				tuser_save	[	241	]	<=	tuser_save	[	240	]	;
				tuser_save	[	242	]	<=	tuser_save	[	241	]	;
				tuser_save	[	243	]	<=	tuser_save	[	242	]	;
				tuser_save	[	244	]	<=	tuser_save	[	243	]	;
				tuser_save	[	245	]	<=	tuser_save	[	244	]	;
				tuser_save	[	246	]	<=	tuser_save	[	245	]	;
				tuser_save	[	247	]	<=	tuser_save	[	246	]	;
				tuser_save	[	248	]	<=	tuser_save	[	247	]	;
				tuser_save	[	249	]	<=	tuser_save	[	248	]	;
				tuser_save	[	250	]	<=	tuser_save	[	249	]	;
				tuser_save	[	251	]	<=	tuser_save	[	250	]	;
				tuser_save	[	252	]	<=	tuser_save	[	251	]	;
				tuser_save	[	253	]	<=	tuser_save	[	252	]	;
				tuser_save	[	254	]	<=	tuser_save	[	253	]	;
				tuser_save	[	255	]	<=	tuser_save	[	254	]	;
					count_packet	<= 2'd0;
					sum_tdata		<=	tdata_save[255];
					sum_tuser		<=	tuser_save[127];
					if(tuser_save[127] == 128'd0)
					begin
						sum_tdata_valid		<=	1'b0;
						sum_tuser_valid		<=	1'b0;
					end
					else
					begin
						sum_tdata_valid		<=	1'b1;
						sum_tuser_valid		<=	1'b1;
					end
				end
			end
		end
		else
		begin
			if(tdata_save[255] == 201'd0)
			begin
				tdata_save	[	0	]	<=	tdata_save	[	0	]	;//stay_no_change
					tdata_save	[	1	]	<=	tdata_save	[	1	]	;
					tdata_save	[	2	]	<=	tdata_save	[	2	]	;
					tdata_save	[	3	]	<=	tdata_save	[	3	]	;
					tdata_save	[	4	]	<=	tdata_save	[	4	]	;
					tdata_save	[	5	]	<=	tdata_save	[	5	]	;
					tdata_save	[	6	]	<=	tdata_save	[	6	]	;
					tdata_save	[	7	]	<=	tdata_save	[	7	]	;
					tdata_save	[	8	]	<=	tdata_save	[	8	]	;
					tdata_save	[	9	]	<=	tdata_save	[	9	]	;
					tdata_save	[	10	]	<=	tdata_save	[	10	]	;
					tdata_save	[	11	]	<=	tdata_save	[	11	]	;
					tdata_save	[	12	]	<=	tdata_save	[	12	]	;
					tdata_save	[	13	]	<=	tdata_save	[	13	]	;
					tdata_save	[	14	]	<=	tdata_save	[	14	]	;
					tdata_save	[	15	]	<=	tdata_save	[	15	]	;
					tdata_save	[	16	]	<=	tdata_save	[	16	]	;
					tdata_save	[	17	]	<=	tdata_save	[	17	]	;
					tdata_save	[	18	]	<=	tdata_save	[	18	]	;
					tdata_save	[	19	]	<=	tdata_save	[	19	]	;
					tdata_save	[	20	]	<=	tdata_save	[	20	]	;
					tdata_save	[	21	]	<=	tdata_save	[	21	]	;
					tdata_save	[	22	]	<=	tdata_save	[	22	]	;
					tdata_save	[	23	]	<=	tdata_save	[	23	]	;
					tdata_save	[	24	]	<=	tdata_save	[	24	]	;
					tdata_save	[	25	]	<=	tdata_save	[	25	]	;
					tdata_save	[	26	]	<=	tdata_save	[	26	]	;
					tdata_save	[	27	]	<=	tdata_save	[	27	]	;
					tdata_save	[	28	]	<=	tdata_save	[	28	]	;
					tdata_save	[	29	]	<=	tdata_save	[	29	]	;
					tdata_save	[	30	]	<=	tdata_save	[	30	]	;
					tdata_save	[	31	]	<=	tdata_save	[	31	]	;
					tdata_save	[	32	]	<=	tdata_save	[	32	]	;
					tdata_save	[	33	]	<=	tdata_save	[	33	]	;
					tdata_save	[	34	]	<=	tdata_save	[	34	]	;
					tdata_save	[	35	]	<=	tdata_save	[	35	]	;
					tdata_save	[	36	]	<=	tdata_save	[	36	]	;
					tdata_save	[	37	]	<=	tdata_save	[	37	]	;
					tdata_save	[	38	]	<=	tdata_save	[	38	]	;
					tdata_save	[	39	]	<=	tdata_save	[	39	]	;
					tdata_save	[	40	]	<=	tdata_save	[	40	]	;
					tdata_save	[	41	]	<=	tdata_save	[	41	]	;
					tdata_save	[	42	]	<=	tdata_save	[	42	]	;
					tdata_save	[	43	]	<=	tdata_save	[	43	]	;
					tdata_save	[	44	]	<=	tdata_save	[	44	]	;
					tdata_save	[	45	]	<=	tdata_save	[	45	]	;
					tdata_save	[	46	]	<=	tdata_save	[	46	]	;
					tdata_save	[	47	]	<=	tdata_save	[	47	]	;
					tdata_save	[	48	]	<=	tdata_save	[	48	]	;
					tdata_save	[	49	]	<=	tdata_save	[	49	]	;
					tdata_save	[	50	]	<=	tdata_save	[	50	]	;
					tdata_save	[	51	]	<=	tdata_save	[	51	]	;
					tdata_save	[	52	]	<=	tdata_save	[	52	]	;
					tdata_save	[	53	]	<=	tdata_save	[	53	]	;
					tdata_save	[	54	]	<=	tdata_save	[	54	]	;
					tdata_save	[	55	]	<=	tdata_save	[	55	]	;
					tdata_save	[	56	]	<=	tdata_save	[	56	]	;
					tdata_save	[	57	]	<=	tdata_save	[	57	]	;
					tdata_save	[	58	]	<=	tdata_save	[	58	]	;
					tdata_save	[	59	]	<=	tdata_save	[	59	]	;
					tdata_save	[	60	]	<=	tdata_save	[	60	]	;
					tdata_save	[	61	]	<=	tdata_save	[	61	]	;
					tdata_save	[	62	]	<=	tdata_save	[	62	]	;
					tdata_save	[	63	]	<=	tdata_save	[	63	]	;
					tdata_save	[	64	]	<=	tdata_save	[	64	]	;
					tdata_save	[	65	]	<=	tdata_save	[	65	]	;
					tdata_save	[	66	]	<=	tdata_save	[	66	]	;
					tdata_save	[	67	]	<=	tdata_save	[	67	]	;
					tdata_save	[	68	]	<=	tdata_save	[	68	]	;
					tdata_save	[	69	]	<=	tdata_save	[	69	]	;
					tdata_save	[	70	]	<=	tdata_save	[	70	]	;
					tdata_save	[	71	]	<=	tdata_save	[	71	]	;
					tdata_save	[	72	]	<=	tdata_save	[	72	]	;
					tdata_save	[	73	]	<=	tdata_save	[	73	]	;
					tdata_save	[	74	]	<=	tdata_save	[	74	]	;
					tdata_save	[	75	]	<=	tdata_save	[	75	]	;
					tdata_save	[	76	]	<=	tdata_save	[	76	]	;
					tdata_save	[	77	]	<=	tdata_save	[	77	]	;
					tdata_save	[	78	]	<=	tdata_save	[	78	]	;
					tdata_save	[	79	]	<=	tdata_save	[	79	]	;
					tdata_save	[	80	]	<=	tdata_save	[	80	]	;
					tdata_save	[	81	]	<=	tdata_save	[	81	]	;
					tdata_save	[	82	]	<=	tdata_save	[	82	]	;
					tdata_save	[	83	]	<=	tdata_save	[	83	]	;
					tdata_save	[	84	]	<=	tdata_save	[	84	]	;
					tdata_save	[	85	]	<=	tdata_save	[	85	]	;
					tdata_save	[	86	]	<=	tdata_save	[	86	]	;
					tdata_save	[	87	]	<=	tdata_save	[	87	]	;
					tdata_save	[	88	]	<=	tdata_save	[	88	]	;
					tdata_save	[	89	]	<=	tdata_save	[	89	]	;
					tdata_save	[	90	]	<=	tdata_save	[	90	]	;
					tdata_save	[	91	]	<=	tdata_save	[	91	]	;
					tdata_save	[	92	]	<=	tdata_save	[	92	]	;
					tdata_save	[	93	]	<=	tdata_save	[	93	]	;
					tdata_save	[	94	]	<=	tdata_save	[	94	]	;
					tdata_save	[	95	]	<=	tdata_save	[	95	]	;
					tdata_save	[	96	]	<=	tdata_save	[	96	]	;
					tdata_save	[	97	]	<=	tdata_save	[	97	]	;
					tdata_save	[	98	]	<=	tdata_save	[	98	]	;
					tdata_save	[	99	]	<=	tdata_save	[	99	]	;
					tdata_save	[	100	]	<=	tdata_save	[	100	]	;
					tdata_save	[	101	]	<=	tdata_save	[	101	]	;
					tdata_save	[	102	]	<=	tdata_save	[	102	]	;
					tdata_save	[	103	]	<=	tdata_save	[	103	]	;
					tdata_save	[	104	]	<=	tdata_save	[	104	]	;
					tdata_save	[	105	]	<=	tdata_save	[	105	]	;
					tdata_save	[	106	]	<=	tdata_save	[	106	]	;
					tdata_save	[	107	]	<=	tdata_save	[	107	]	;
					tdata_save	[	108	]	<=	tdata_save	[	108	]	;
					tdata_save	[	109	]	<=	tdata_save	[	109	]	;
					tdata_save	[	110	]	<=	tdata_save	[	110	]	;
					tdata_save	[	111	]	<=	tdata_save	[	111	]	;
					tdata_save	[	112	]	<=	tdata_save	[	112	]	;
					tdata_save	[	113	]	<=	tdata_save	[	113	]	;
					tdata_save	[	114	]	<=	tdata_save	[	114	]	;
					tdata_save	[	115	]	<=	tdata_save	[	115	]	;
					tdata_save	[	116	]	<=	tdata_save	[	116	]	;
					tdata_save	[	117	]	<=	tdata_save	[	117	]	;
					tdata_save	[	118	]	<=	tdata_save	[	118	]	;
					tdata_save	[	119	]	<=	tdata_save	[	119	]	;
					tdata_save	[	120	]	<=	tdata_save	[	120	]	;
					tdata_save	[	121	]	<=	tdata_save	[	121	]	;
					tdata_save	[	122	]	<=	tdata_save	[	122	]	;
					tdata_save	[	123	]	<=	tdata_save	[	123	]	;
					tdata_save	[	124	]	<=	tdata_save	[	124	]	;
					tdata_save	[	125	]	<=	tdata_save	[	125	]	;
					tdata_save	[	126	]	<=	tdata_save	[	126	]	;
					tdata_save	[	127	]	<=	tdata_save	[	127	]	;
					tdata_save	[	128	]	<=	tdata_save	[	128	]	;
					tdata_save	[	129	]	<=	tdata_save	[	129	]	;
					tdata_save	[	130	]	<=	tdata_save	[	130	]	;
					tdata_save	[	131	]	<=	tdata_save	[	131	]	;
					tdata_save	[	132	]	<=	tdata_save	[	132	]	;
					tdata_save	[	133	]	<=	tdata_save	[	133	]	;
					tdata_save	[	134	]	<=	tdata_save	[	134	]	;
					tdata_save	[	135	]	<=	tdata_save	[	135	]	;
					tdata_save	[	136	]	<=	tdata_save	[	136	]	;
					tdata_save	[	137	]	<=	tdata_save	[	137	]	;
					tdata_save	[	138	]	<=	tdata_save	[	138	]	;
					tdata_save	[	139	]	<=	tdata_save	[	139	]	;
					tdata_save	[	140	]	<=	tdata_save	[	140	]	;
					tdata_save	[	141	]	<=	tdata_save	[	141	]	;
					tdata_save	[	142	]	<=	tdata_save	[	142	]	;
					tdata_save	[	143	]	<=	tdata_save	[	143	]	;
					tdata_save	[	144	]	<=	tdata_save	[	144	]	;
					tdata_save	[	145	]	<=	tdata_save	[	145	]	;
					tdata_save	[	146	]	<=	tdata_save	[	146	]	;
					tdata_save	[	147	]	<=	tdata_save	[	147	]	;
					tdata_save	[	148	]	<=	tdata_save	[	148	]	;
					tdata_save	[	149	]	<=	tdata_save	[	149	]	;
					tdata_save	[	150	]	<=	tdata_save	[	150	]	;
					tdata_save	[	151	]	<=	tdata_save	[	151	]	;
					tdata_save	[	152	]	<=	tdata_save	[	152	]	;
					tdata_save	[	153	]	<=	tdata_save	[	153	]	;
					tdata_save	[	154	]	<=	tdata_save	[	154	]	;
					tdata_save	[	155	]	<=	tdata_save	[	155	]	;
					tdata_save	[	156	]	<=	tdata_save	[	156	]	;
					tdata_save	[	157	]	<=	tdata_save	[	157	]	;
					tdata_save	[	158	]	<=	tdata_save	[	158	]	;
					tdata_save	[	159	]	<=	tdata_save	[	159	]	;
					tdata_save	[	160	]	<=	tdata_save	[	160	]	;
					tdata_save	[	161	]	<=	tdata_save	[	161	]	;
					tdata_save	[	162	]	<=	tdata_save	[	162	]	;
					tdata_save	[	163	]	<=	tdata_save	[	163	]	;
					tdata_save	[	164	]	<=	tdata_save	[	164	]	;
					tdata_save	[	165	]	<=	tdata_save	[	165	]	;
					tdata_save	[	166	]	<=	tdata_save	[	166	]	;
					tdata_save	[	167	]	<=	tdata_save	[	167	]	;
					tdata_save	[	168	]	<=	tdata_save	[	168	]	;
					tdata_save	[	169	]	<=	tdata_save	[	169	]	;
					tdata_save	[	170	]	<=	tdata_save	[	170	]	;
					tdata_save	[	171	]	<=	tdata_save	[	171	]	;
					tdata_save	[	172	]	<=	tdata_save	[	172	]	;
					tdata_save	[	173	]	<=	tdata_save	[	173	]	;
					tdata_save	[	174	]	<=	tdata_save	[	174	]	;
					tdata_save	[	175	]	<=	tdata_save	[	175	]	;
					tdata_save	[	176	]	<=	tdata_save	[	176	]	;
					tdata_save	[	177	]	<=	tdata_save	[	177	]	;
					tdata_save	[	178	]	<=	tdata_save	[	178	]	;
					tdata_save	[	179	]	<=	tdata_save	[	179	]	;
					tdata_save	[	180	]	<=	tdata_save	[	180	]	;
					tdata_save	[	181	]	<=	tdata_save	[	181	]	;
					tdata_save	[	182	]	<=	tdata_save	[	182	]	;
					tdata_save	[	183	]	<=	tdata_save	[	183	]	;
					tdata_save	[	184	]	<=	tdata_save	[	184	]	;
					tdata_save	[	185	]	<=	tdata_save	[	185	]	;
					tdata_save	[	186	]	<=	tdata_save	[	186	]	;
					tdata_save	[	187	]	<=	tdata_save	[	187	]	;
					tdata_save	[	188	]	<=	tdata_save	[	188	]	;
					tdata_save	[	189	]	<=	tdata_save	[	189	]	;
					tdata_save	[	190	]	<=	tdata_save	[	190	]	;
					tdata_save	[	191	]	<=	tdata_save	[	191	]	;
					tdata_save	[	192	]	<=	tdata_save	[	192	]	;
					tdata_save	[	193	]	<=	tdata_save	[	193	]	;
					tdata_save	[	194	]	<=	tdata_save	[	194	]	;
					tdata_save	[	195	]	<=	tdata_save	[	195	]	;
					tdata_save	[	196	]	<=	tdata_save	[	196	]	;
					tdata_save	[	197	]	<=	tdata_save	[	197	]	;
					tdata_save	[	198	]	<=	tdata_save	[	198	]	;
					tdata_save	[	199	]	<=	tdata_save	[	199	]	;
					tdata_save	[	200	]	<=	tdata_save	[	200	]	;
					tdata_save	[	201	]	<=	tdata_save	[	201	]	;
					tdata_save	[	202	]	<=	tdata_save	[	202	]	;
					tdata_save	[	203	]	<=	tdata_save	[	203	]	;
					tdata_save	[	204	]	<=	tdata_save	[	204	]	;
					tdata_save	[	205	]	<=	tdata_save	[	205	]	;
					tdata_save	[	206	]	<=	tdata_save	[	206	]	;
					tdata_save	[	207	]	<=	tdata_save	[	207	]	;
					tdata_save	[	208	]	<=	tdata_save	[	208	]	;
					tdata_save	[	209	]	<=	tdata_save	[	209	]	;
					tdata_save	[	210	]	<=	tdata_save	[	210	]	;
					tdata_save	[	211	]	<=	tdata_save	[	211	]	;
					tdata_save	[	212	]	<=	tdata_save	[	212	]	;
					tdata_save	[	213	]	<=	tdata_save	[	213	]	;
					tdata_save	[	214	]	<=	tdata_save	[	214	]	;
					tdata_save	[	215	]	<=	tdata_save	[	215	]	;
					tdata_save	[	216	]	<=	tdata_save	[	216	]	;
					tdata_save	[	217	]	<=	tdata_save	[	217	]	;
					tdata_save	[	218	]	<=	tdata_save	[	218	]	;
					tdata_save	[	219	]	<=	tdata_save	[	219	]	;
					tdata_save	[	220	]	<=	tdata_save	[	220	]	;
					tdata_save	[	221	]	<=	tdata_save	[	221	]	;
					tdata_save	[	222	]	<=	tdata_save	[	222	]	;
					tdata_save	[	223	]	<=	tdata_save	[	223	]	;
					tdata_save	[	224	]	<=	tdata_save	[	224	]	;
					tdata_save	[	225	]	<=	tdata_save	[	225	]	;
					tdata_save	[	226	]	<=	tdata_save	[	226	]	;
					tdata_save	[	227	]	<=	tdata_save	[	227	]	;
					tdata_save	[	228	]	<=	tdata_save	[	228	]	;
					tdata_save	[	229	]	<=	tdata_save	[	229	]	;
					tdata_save	[	230	]	<=	tdata_save	[	230	]	;
					tdata_save	[	231	]	<=	tdata_save	[	231	]	;
					tdata_save	[	232	]	<=	tdata_save	[	232	]	;
					tdata_save	[	233	]	<=	tdata_save	[	233	]	;
					tdata_save	[	234	]	<=	tdata_save	[	234	]	;
					tdata_save	[	235	]	<=	tdata_save	[	235	]	;
					tdata_save	[	236	]	<=	tdata_save	[	236	]	;
					tdata_save	[	237	]	<=	tdata_save	[	237	]	;
					tdata_save	[	238	]	<=	tdata_save	[	238	]	;
					tdata_save	[	239	]	<=	tdata_save	[	239	]	;
					tdata_save	[	240	]	<=	tdata_save	[	240	]	;
					tdata_save	[	241	]	<=	tdata_save	[	241	]	;
					tdata_save	[	242	]	<=	tdata_save	[	242	]	;
					tdata_save	[	243	]	<=	tdata_save	[	243	]	;
					tdata_save	[	244	]	<=	tdata_save	[	244	]	;
					tdata_save	[	245	]	<=	tdata_save	[	245	]	;
					tdata_save	[	246	]	<=	tdata_save	[	246	]	;
					tdata_save	[	247	]	<=	tdata_save	[	247	]	;
					tdata_save	[	248	]	<=	tdata_save	[	248	]	;
					tdata_save	[	249	]	<=	tdata_save	[	249	]	;
					tdata_save	[	250	]	<=	tdata_save	[	250	]	;
					tdata_save	[	251	]	<=	tdata_save	[	251	]	;
					tdata_save	[	252	]	<=	tdata_save	[	252	]	;
					tdata_save	[	253	]	<=	tdata_save	[	253	]	;
					tdata_save	[	254	]	<=	tdata_save	[	254	]	;
					tdata_save	[	255	]	<=	tdata_save	[	255	]	;
				tuser_save	[	0	]	<=	tuser_save	[	0	]	;
				tuser_save	[	1	]	<=	tuser_save	[	1	]	;
				tuser_save	[	2	]	<=	tuser_save	[	2	]	;
				tuser_save	[	3	]	<=	tuser_save	[	3	]	;
				tuser_save	[	4	]	<=	tuser_save	[	4	]	;
				tuser_save	[	5	]	<=	tuser_save	[	5	]	;
				tuser_save	[	6	]	<=	tuser_save	[	6	]	;
				tuser_save	[	7	]	<=	tuser_save	[	7	]	;
				tuser_save	[	8	]	<=	tuser_save	[	8	]	;
				tuser_save	[	9	]	<=	tuser_save	[	9	]	;
				tuser_save	[	10	]	<=	tuser_save	[	10	]	;
				tuser_save	[	11	]	<=	tuser_save	[	11	]	;
				tuser_save	[	12	]	<=	tuser_save	[	12	]	;
				tuser_save	[	13	]	<=	tuser_save	[	13	]	;
				tuser_save	[	14	]	<=	tuser_save	[	14	]	;
				tuser_save	[	15	]	<=	tuser_save	[	15	]	;
				tuser_save	[	16	]	<=	tuser_save	[	16	]	;
				tuser_save	[	17	]	<=	tuser_save	[	17	]	;
				tuser_save	[	18	]	<=	tuser_save	[	18	]	;
				tuser_save	[	19	]	<=	tuser_save	[	19	]	;
				tuser_save	[	20	]	<=	tuser_save	[	20	]	;
				tuser_save	[	21	]	<=	tuser_save	[	21	]	;
				tuser_save	[	22	]	<=	tuser_save	[	22	]	;
				tuser_save	[	23	]	<=	tuser_save	[	23	]	;
				tuser_save	[	24	]	<=	tuser_save	[	24	]	;
				tuser_save	[	25	]	<=	tuser_save	[	25	]	;
				tuser_save	[	26	]	<=	tuser_save	[	26	]	;
				tuser_save	[	27	]	<=	tuser_save	[	27	]	;
				tuser_save	[	28	]	<=	tuser_save	[	28	]	;
				tuser_save	[	29	]	<=	tuser_save	[	29	]	;
				tuser_save	[	30	]	<=	tuser_save	[	30	]	;
				tuser_save	[	31	]	<=	tuser_save	[	31	]	;
				tuser_save	[	32	]	<=	tuser_save	[	32	]	;
				tuser_save	[	33	]	<=	tuser_save	[	33	]	;
				tuser_save	[	34	]	<=	tuser_save	[	34	]	;
				tuser_save	[	35	]	<=	tuser_save	[	35	]	;
				tuser_save	[	36	]	<=	tuser_save	[	36	]	;
				tuser_save	[	37	]	<=	tuser_save	[	37	]	;
				tuser_save	[	38	]	<=	tuser_save	[	38	]	;
				tuser_save	[	39	]	<=	tuser_save	[	39	]	;
				tuser_save	[	40	]	<=	tuser_save	[	40	]	;
				tuser_save	[	41	]	<=	tuser_save	[	41	]	;
				tuser_save	[	42	]	<=	tuser_save	[	42	]	;
				tuser_save	[	43	]	<=	tuser_save	[	43	]	;
				tuser_save	[	44	]	<=	tuser_save	[	44	]	;
				tuser_save	[	45	]	<=	tuser_save	[	45	]	;
				tuser_save	[	46	]	<=	tuser_save	[	46	]	;
				tuser_save	[	47	]	<=	tuser_save	[	47	]	;
				tuser_save	[	48	]	<=	tuser_save	[	48	]	;
				tuser_save	[	49	]	<=	tuser_save	[	49	]	;
				tuser_save	[	50	]	<=	tuser_save	[	50	]	;
				tuser_save	[	51	]	<=	tuser_save	[	51	]	;
				tuser_save	[	52	]	<=	tuser_save	[	52	]	;
				tuser_save	[	53	]	<=	tuser_save	[	53	]	;
				tuser_save	[	54	]	<=	tuser_save	[	54	]	;
				tuser_save	[	55	]	<=	tuser_save	[	55	]	;
				tuser_save	[	56	]	<=	tuser_save	[	56	]	;
				tuser_save	[	57	]	<=	tuser_save	[	57	]	;
				tuser_save	[	58	]	<=	tuser_save	[	58	]	;
				tuser_save	[	59	]	<=	tuser_save	[	59	]	;
				tuser_save	[	60	]	<=	tuser_save	[	60	]	;
				tuser_save	[	61	]	<=	tuser_save	[	61	]	;
				tuser_save	[	62	]	<=	tuser_save	[	62	]	;
				tuser_save	[	63	]	<=	tuser_save	[	63	]	;
				tuser_save	[	64	]	<=	tuser_save	[	64	]	;
				tuser_save	[	65	]	<=	tuser_save	[	65	]	;
				tuser_save	[	66	]	<=	tuser_save	[	66	]	;
				tuser_save	[	67	]	<=	tuser_save	[	67	]	;
				tuser_save	[	68	]	<=	tuser_save	[	68	]	;
				tuser_save	[	69	]	<=	tuser_save	[	69	]	;
				tuser_save	[	70	]	<=	tuser_save	[	70	]	;
				tuser_save	[	71	]	<=	tuser_save	[	71	]	;
				tuser_save	[	72	]	<=	tuser_save	[	72	]	;
				tuser_save	[	73	]	<=	tuser_save	[	73	]	;
				tuser_save	[	74	]	<=	tuser_save	[	74	]	;
				tuser_save	[	75	]	<=	tuser_save	[	75	]	;
				tuser_save	[	76	]	<=	tuser_save	[	76	]	;
				tuser_save	[	77	]	<=	tuser_save	[	77	]	;
				tuser_save	[	78	]	<=	tuser_save	[	78	]	;
				tuser_save	[	79	]	<=	tuser_save	[	79	]	;
				tuser_save	[	80	]	<=	tuser_save	[	80	]	;
				tuser_save	[	81	]	<=	tuser_save	[	81	]	;
				tuser_save	[	82	]	<=	tuser_save	[	82	]	;
				tuser_save	[	83	]	<=	tuser_save	[	83	]	;
				tuser_save	[	84	]	<=	tuser_save	[	84	]	;
				tuser_save	[	85	]	<=	tuser_save	[	85	]	;
				tuser_save	[	86	]	<=	tuser_save	[	86	]	;
				tuser_save	[	87	]	<=	tuser_save	[	87	]	;
				tuser_save	[	88	]	<=	tuser_save	[	88	]	;
				tuser_save	[	89	]	<=	tuser_save	[	89	]	;
				tuser_save	[	90	]	<=	tuser_save	[	90	]	;
				tuser_save	[	91	]	<=	tuser_save	[	91	]	;
				tuser_save	[	92	]	<=	tuser_save	[	92	]	;
				tuser_save	[	93	]	<=	tuser_save	[	93	]	;
				tuser_save	[	94	]	<=	tuser_save	[	94	]	;
				tuser_save	[	95	]	<=	tuser_save	[	95	]	;
				tuser_save	[	96	]	<=	tuser_save	[	96	]	;
				tuser_save	[	97	]	<=	tuser_save	[	97	]	;
				tuser_save	[	98	]	<=	tuser_save	[	98	]	;
				tuser_save	[	99	]	<=	tuser_save	[	99	]	;
				tuser_save	[	100	]	<=	tuser_save	[	100	]	;
				tuser_save	[	101	]	<=	tuser_save	[	101	]	;
				tuser_save	[	102	]	<=	tuser_save	[	102	]	;
				tuser_save	[	103	]	<=	tuser_save	[	103	]	;
				tuser_save	[	104	]	<=	tuser_save	[	104	]	;
				tuser_save	[	105	]	<=	tuser_save	[	105	]	;
				tuser_save	[	106	]	<=	tuser_save	[	106	]	;
				tuser_save	[	107	]	<=	tuser_save	[	107	]	;
				tuser_save	[	108	]	<=	tuser_save	[	108	]	;
				tuser_save	[	109	]	<=	tuser_save	[	109	]	;
				tuser_save	[	110	]	<=	tuser_save	[	110	]	;
				tuser_save	[	111	]	<=	tuser_save	[	111	]	;
				tuser_save	[	112	]	<=	tuser_save	[	112	]	;
				tuser_save	[	113	]	<=	tuser_save	[	113	]	;
				tuser_save	[	114	]	<=	tuser_save	[	114	]	;
				tuser_save	[	115	]	<=	tuser_save	[	115	]	;
				tuser_save	[	116	]	<=	tuser_save	[	116	]	;
				tuser_save	[	117	]	<=	tuser_save	[	117	]	;
				tuser_save	[	118	]	<=	tuser_save	[	118	]	;
				tuser_save	[	119	]	<=	tuser_save	[	119	]	;
				tuser_save	[	120	]	<=	tuser_save	[	120	]	;
				tuser_save	[	121	]	<=	tuser_save	[	121	]	;
				tuser_save	[	122	]	<=	tuser_save	[	122	]	;
				tuser_save	[	123	]	<=	tuser_save	[	123	]	;
				tuser_save	[	124	]	<=	tuser_save	[	124	]	;
				tuser_save	[	125	]	<=	tuser_save	[	125	]	;
				tuser_save	[	126	]	<=	tuser_save	[	126	]	;
				tuser_save	[	127	]	<=	tuser_save	[	127	]	;
				tuser_save	[	128	]	<=	tuser_save	[	128	]	;
				tuser_save	[	129	]	<=	tuser_save	[	129	]	;
				tuser_save	[	130	]	<=	tuser_save	[	130	]	;
				tuser_save	[	131	]	<=	tuser_save	[	131	]	;
				tuser_save	[	132	]	<=	tuser_save	[	132	]	;
				tuser_save	[	133	]	<=	tuser_save	[	133	]	;
				tuser_save	[	134	]	<=	tuser_save	[	134	]	;
				tuser_save	[	135	]	<=	tuser_save	[	135	]	;
				tuser_save	[	136	]	<=	tuser_save	[	136	]	;
				tuser_save	[	137	]	<=	tuser_save	[	137	]	;
				tuser_save	[	138	]	<=	tuser_save	[	138	]	;
				tuser_save	[	139	]	<=	tuser_save	[	139	]	;
				tuser_save	[	140	]	<=	tuser_save	[	140	]	;
				tuser_save	[	141	]	<=	tuser_save	[	141	]	;
				tuser_save	[	142	]	<=	tuser_save	[	142	]	;
				tuser_save	[	143	]	<=	tuser_save	[	143	]	;
				tuser_save	[	144	]	<=	tuser_save	[	144	]	;
				tuser_save	[	145	]	<=	tuser_save	[	145	]	;
				tuser_save	[	146	]	<=	tuser_save	[	146	]	;
				tuser_save	[	147	]	<=	tuser_save	[	147	]	;
				tuser_save	[	148	]	<=	tuser_save	[	148	]	;
				tuser_save	[	149	]	<=	tuser_save	[	149	]	;
				tuser_save	[	150	]	<=	tuser_save	[	150	]	;
				tuser_save	[	151	]	<=	tuser_save	[	151	]	;
				tuser_save	[	152	]	<=	tuser_save	[	152	]	;
				tuser_save	[	153	]	<=	tuser_save	[	153	]	;
				tuser_save	[	154	]	<=	tuser_save	[	154	]	;
				tuser_save	[	155	]	<=	tuser_save	[	155	]	;
				tuser_save	[	156	]	<=	tuser_save	[	156	]	;
				tuser_save	[	157	]	<=	tuser_save	[	157	]	;
				tuser_save	[	158	]	<=	tuser_save	[	158	]	;
				tuser_save	[	159	]	<=	tuser_save	[	159	]	;
				tuser_save	[	160	]	<=	tuser_save	[	160	]	;
				tuser_save	[	161	]	<=	tuser_save	[	161	]	;
				tuser_save	[	162	]	<=	tuser_save	[	162	]	;
				tuser_save	[	163	]	<=	tuser_save	[	163	]	;
				tuser_save	[	164	]	<=	tuser_save	[	164	]	;
				tuser_save	[	165	]	<=	tuser_save	[	165	]	;
				tuser_save	[	166	]	<=	tuser_save	[	166	]	;
				tuser_save	[	167	]	<=	tuser_save	[	167	]	;
				tuser_save	[	168	]	<=	tuser_save	[	168	]	;
				tuser_save	[	169	]	<=	tuser_save	[	169	]	;
				tuser_save	[	170	]	<=	tuser_save	[	170	]	;
				tuser_save	[	171	]	<=	tuser_save	[	171	]	;
				tuser_save	[	172	]	<=	tuser_save	[	172	]	;
				tuser_save	[	173	]	<=	tuser_save	[	173	]	;
				tuser_save	[	174	]	<=	tuser_save	[	174	]	;
				tuser_save	[	175	]	<=	tuser_save	[	175	]	;
				tuser_save	[	176	]	<=	tuser_save	[	176	]	;
				tuser_save	[	177	]	<=	tuser_save	[	177	]	;
				tuser_save	[	178	]	<=	tuser_save	[	178	]	;
				tuser_save	[	179	]	<=	tuser_save	[	179	]	;
				tuser_save	[	180	]	<=	tuser_save	[	180	]	;
				tuser_save	[	181	]	<=	tuser_save	[	181	]	;
				tuser_save	[	182	]	<=	tuser_save	[	182	]	;
				tuser_save	[	183	]	<=	tuser_save	[	183	]	;
				tuser_save	[	184	]	<=	tuser_save	[	184	]	;
				tuser_save	[	185	]	<=	tuser_save	[	185	]	;
				tuser_save	[	186	]	<=	tuser_save	[	186	]	;
				tuser_save	[	187	]	<=	tuser_save	[	187	]	;
				tuser_save	[	188	]	<=	tuser_save	[	188	]	;
				tuser_save	[	189	]	<=	tuser_save	[	189	]	;
				tuser_save	[	190	]	<=	tuser_save	[	190	]	;
				tuser_save	[	191	]	<=	tuser_save	[	191	]	;
				tuser_save	[	192	]	<=	tuser_save	[	192	]	;
				tuser_save	[	193	]	<=	tuser_save	[	193	]	;
				tuser_save	[	194	]	<=	tuser_save	[	194	]	;
				tuser_save	[	195	]	<=	tuser_save	[	195	]	;
				tuser_save	[	196	]	<=	tuser_save	[	196	]	;
				tuser_save	[	197	]	<=	tuser_save	[	197	]	;
				tuser_save	[	198	]	<=	tuser_save	[	198	]	;
				tuser_save	[	199	]	<=	tuser_save	[	199	]	;
				tuser_save	[	200	]	<=	tuser_save	[	200	]	;
				tuser_save	[	201	]	<=	tuser_save	[	201	]	;
				tuser_save	[	202	]	<=	tuser_save	[	202	]	;
				tuser_save	[	203	]	<=	tuser_save	[	203	]	;
				tuser_save	[	204	]	<=	tuser_save	[	204	]	;
				tuser_save	[	205	]	<=	tuser_save	[	205	]	;
				tuser_save	[	206	]	<=	tuser_save	[	206	]	;
				tuser_save	[	207	]	<=	tuser_save	[	207	]	;
				tuser_save	[	208	]	<=	tuser_save	[	208	]	;
				tuser_save	[	209	]	<=	tuser_save	[	209	]	;
				tuser_save	[	210	]	<=	tuser_save	[	210	]	;
				tuser_save	[	211	]	<=	tuser_save	[	211	]	;
				tuser_save	[	212	]	<=	tuser_save	[	212	]	;
				tuser_save	[	213	]	<=	tuser_save	[	213	]	;
				tuser_save	[	214	]	<=	tuser_save	[	214	]	;
				tuser_save	[	215	]	<=	tuser_save	[	215	]	;
				tuser_save	[	216	]	<=	tuser_save	[	216	]	;
				tuser_save	[	217	]	<=	tuser_save	[	217	]	;
				tuser_save	[	218	]	<=	tuser_save	[	218	]	;
				tuser_save	[	219	]	<=	tuser_save	[	219	]	;
				tuser_save	[	220	]	<=	tuser_save	[	220	]	;
				tuser_save	[	221	]	<=	tuser_save	[	221	]	;
				tuser_save	[	222	]	<=	tuser_save	[	222	]	;
				tuser_save	[	223	]	<=	tuser_save	[	223	]	;
				tuser_save	[	224	]	<=	tuser_save	[	224	]	;
				tuser_save	[	225	]	<=	tuser_save	[	225	]	;
				tuser_save	[	226	]	<=	tuser_save	[	226	]	;
				tuser_save	[	227	]	<=	tuser_save	[	227	]	;
				tuser_save	[	228	]	<=	tuser_save	[	228	]	;
				tuser_save	[	229	]	<=	tuser_save	[	229	]	;
				tuser_save	[	230	]	<=	tuser_save	[	230	]	;
				tuser_save	[	231	]	<=	tuser_save	[	231	]	;
				tuser_save	[	232	]	<=	tuser_save	[	232	]	;
				tuser_save	[	233	]	<=	tuser_save	[	233	]	;
				tuser_save	[	234	]	<=	tuser_save	[	234	]	;
				tuser_save	[	235	]	<=	tuser_save	[	235	]	;
				tuser_save	[	236	]	<=	tuser_save	[	236	]	;
				tuser_save	[	237	]	<=	tuser_save	[	237	]	;
				tuser_save	[	238	]	<=	tuser_save	[	238	]	;
				tuser_save	[	239	]	<=	tuser_save	[	239	]	;
				tuser_save	[	240	]	<=	tuser_save	[	240	]	;
				tuser_save	[	241	]	<=	tuser_save	[	241	]	;
				tuser_save	[	242	]	<=	tuser_save	[	242	]	;
				tuser_save	[	243	]	<=	tuser_save	[	243	]	;
				tuser_save	[	244	]	<=	tuser_save	[	244	]	;
				tuser_save	[	245	]	<=	tuser_save	[	245	]	;
				tuser_save	[	246	]	<=	tuser_save	[	246	]	;
				tuser_save	[	247	]	<=	tuser_save	[	247	]	;
				tuser_save	[	248	]	<=	tuser_save	[	248	]	;
				tuser_save	[	249	]	<=	tuser_save	[	249	]	;
				tuser_save	[	250	]	<=	tuser_save	[	250	]	;
				tuser_save	[	251	]	<=	tuser_save	[	251	]	;
				tuser_save	[	252	]	<=	tuser_save	[	252	]	;
				tuser_save	[	253	]	<=	tuser_save	[	253	]	;
				tuser_save	[	254	]	<=	tuser_save	[	254	]	;
				tuser_save	[	255	]	<=	tuser_save	[	255	]	;
				if(count_packet == 2'd2)
					begin
						count_packet <= 2'd0;
					end
					else
					begin
						count_packet	<= count_packet;
					end
				sum_tdata		<=	201'd0;
				sum_tuser		<=	128'd0;
				sum_tdata_valid		<=	1'b0;
				sum_tuser_valid		<=	1'b0;
			end
			else
			begin
				tdata_save	[	0	]	<=	axififo_din;	//shift			
					tdata_save	[	1	]	<=	tdata_save	[	0	]	;
					tdata_save	[	2	]	<=	tdata_save	[	1	]	;
					tdata_save	[	3	]	<=	tdata_save	[	2	]	;
					tdata_save	[	4	]	<=	tdata_save	[	3	]	;
					tdata_save	[	5	]	<=	tdata_save	[	4	]	;
					tdata_save	[	6	]	<=	tdata_save	[	5	]	;
					tdata_save	[	7	]	<=	tdata_save	[	6	]	;
					tdata_save	[	8	]	<=	tdata_save	[	7	]	;
					tdata_save	[	9	]	<=	tdata_save	[	8	]	;
					tdata_save	[	10	]	<=	tdata_save	[	9	]	;
					tdata_save	[	11	]	<=	tdata_save	[	10	]	;
					tdata_save	[	12	]	<=	tdata_save	[	11	]	;
					tdata_save	[	13	]	<=	tdata_save	[	12	]	;
					tdata_save	[	14	]	<=	tdata_save	[	13	]	;
					tdata_save	[	15	]	<=	tdata_save	[	14	]	;
					tdata_save	[	16	]	<=	tdata_save	[	15	]	;
					tdata_save	[	17	]	<=	tdata_save	[	16	]	;
					tdata_save	[	18	]	<=	tdata_save	[	17	]	;
					tdata_save	[	19	]	<=	tdata_save	[	18	]	;
					tdata_save	[	20	]	<=	tdata_save	[	19	]	;
					tdata_save	[	21	]	<=	tdata_save	[	20	]	;
					tdata_save	[	22	]	<=	tdata_save	[	21	]	;
					tdata_save	[	23	]	<=	tdata_save	[	22	]	;
					tdata_save	[	24	]	<=	tdata_save	[	23	]	;
					tdata_save	[	25	]	<=	tdata_save	[	24	]	;
					tdata_save	[	26	]	<=	tdata_save	[	25	]	;
					tdata_save	[	27	]	<=	tdata_save	[	26	]	;
					tdata_save	[	28	]	<=	tdata_save	[	27	]	;
					tdata_save	[	29	]	<=	tdata_save	[	28	]	;
					tdata_save	[	30	]	<=	tdata_save	[	29	]	;
					tdata_save	[	31	]	<=	tdata_save	[	30	]	;
					tdata_save	[	32	]	<=	tdata_save	[	31	]	;
					tdata_save	[	33	]	<=	tdata_save	[	32	]	;
					tdata_save	[	34	]	<=	tdata_save	[	33	]	;
					tdata_save	[	35	]	<=	tdata_save	[	34	]	;
					tdata_save	[	36	]	<=	tdata_save	[	35	]	;
					tdata_save	[	37	]	<=	tdata_save	[	36	]	;
					tdata_save	[	38	]	<=	tdata_save	[	37	]	;
					tdata_save	[	39	]	<=	tdata_save	[	38	]	;
					tdata_save	[	40	]	<=	tdata_save	[	39	]	;
					tdata_save	[	41	]	<=	tdata_save	[	40	]	;
					tdata_save	[	42	]	<=	tdata_save	[	41	]	;
					tdata_save	[	43	]	<=	tdata_save	[	42	]	;
					tdata_save	[	44	]	<=	tdata_save	[	43	]	;
					tdata_save	[	45	]	<=	tdata_save	[	44	]	;
					tdata_save	[	46	]	<=	tdata_save	[	45	]	;
					tdata_save	[	47	]	<=	tdata_save	[	46	]	;
					tdata_save	[	48	]	<=	tdata_save	[	47	]	;
					tdata_save	[	49	]	<=	tdata_save	[	48	]	;
					tdata_save	[	50	]	<=	tdata_save	[	49	]	;
					tdata_save	[	51	]	<=	tdata_save	[	50	]	;
					tdata_save	[	52	]	<=	tdata_save	[	51	]	;
					tdata_save	[	53	]	<=	tdata_save	[	52	]	;
					tdata_save	[	54	]	<=	tdata_save	[	53	]	;
					tdata_save	[	55	]	<=	tdata_save	[	54	]	;
					tdata_save	[	56	]	<=	tdata_save	[	55	]	;
					tdata_save	[	57	]	<=	tdata_save	[	56	]	;
					tdata_save	[	58	]	<=	tdata_save	[	57	]	;
					tdata_save	[	59	]	<=	tdata_save	[	58	]	;
					tdata_save	[	60	]	<=	tdata_save	[	59	]	;
					tdata_save	[	61	]	<=	tdata_save	[	60	]	;
					tdata_save	[	62	]	<=	tdata_save	[	61	]	;
					tdata_save	[	63	]	<=	tdata_save	[	62	]	;
					tdata_save	[	64	]	<=	tdata_save	[	63	]	;
					tdata_save	[	65	]	<=	tdata_save	[	64	]	;
					tdata_save	[	66	]	<=	tdata_save	[	65	]	;
					tdata_save	[	67	]	<=	tdata_save	[	66	]	;
					tdata_save	[	68	]	<=	tdata_save	[	67	]	;
					tdata_save	[	69	]	<=	tdata_save	[	68	]	;
					tdata_save	[	70	]	<=	tdata_save	[	69	]	;
					tdata_save	[	71	]	<=	tdata_save	[	70	]	;
					tdata_save	[	72	]	<=	tdata_save	[	71	]	;
					tdata_save	[	73	]	<=	tdata_save	[	72	]	;
					tdata_save	[	74	]	<=	tdata_save	[	73	]	;
					tdata_save	[	75	]	<=	tdata_save	[	74	]	;
					tdata_save	[	76	]	<=	tdata_save	[	75	]	;
					tdata_save	[	77	]	<=	tdata_save	[	76	]	;
					tdata_save	[	78	]	<=	tdata_save	[	77	]	;
					tdata_save	[	79	]	<=	tdata_save	[	78	]	;
					tdata_save	[	80	]	<=	tdata_save	[	79	]	;
					tdata_save	[	81	]	<=	tdata_save	[	80	]	;
					tdata_save	[	82	]	<=	tdata_save	[	81	]	;
					tdata_save	[	83	]	<=	tdata_save	[	82	]	;
					tdata_save	[	84	]	<=	tdata_save	[	83	]	;
					tdata_save	[	85	]	<=	tdata_save	[	84	]	;
					tdata_save	[	86	]	<=	tdata_save	[	85	]	;
					tdata_save	[	87	]	<=	tdata_save	[	86	]	;
					tdata_save	[	88	]	<=	tdata_save	[	87	]	;
					tdata_save	[	89	]	<=	tdata_save	[	88	]	;
					tdata_save	[	90	]	<=	tdata_save	[	89	]	;
					tdata_save	[	91	]	<=	tdata_save	[	90	]	;
					tdata_save	[	92	]	<=	tdata_save	[	91	]	;
					tdata_save	[	93	]	<=	tdata_save	[	92	]	;
					tdata_save	[	94	]	<=	tdata_save	[	93	]	;
					tdata_save	[	95	]	<=	tdata_save	[	94	]	;
					tdata_save	[	96	]	<=	tdata_save	[	95	]	;
					tdata_save	[	97	]	<=	tdata_save	[	96	]	;
					tdata_save	[	98	]	<=	tdata_save	[	97	]	;
					tdata_save	[	99	]	<=	tdata_save	[	98	]	;
					tdata_save	[	100	]	<=	tdata_save	[	99	]	;
					tdata_save	[	101	]	<=	tdata_save	[	100	]	;
					tdata_save	[	102	]	<=	tdata_save	[	101	]	;
					tdata_save	[	103	]	<=	tdata_save	[	102	]	;
					tdata_save	[	104	]	<=	tdata_save	[	103	]	;
					tdata_save	[	105	]	<=	tdata_save	[	104	]	;
					tdata_save	[	106	]	<=	tdata_save	[	105	]	;
					tdata_save	[	107	]	<=	tdata_save	[	106	]	;
					tdata_save	[	108	]	<=	tdata_save	[	107	]	;
					tdata_save	[	109	]	<=	tdata_save	[	108	]	;
					tdata_save	[	110	]	<=	tdata_save	[	109	]	;
					tdata_save	[	111	]	<=	tdata_save	[	110	]	;
					tdata_save	[	112	]	<=	tdata_save	[	111	]	;
					tdata_save	[	113	]	<=	tdata_save	[	112	]	;
					tdata_save	[	114	]	<=	tdata_save	[	113	]	;
					tdata_save	[	115	]	<=	tdata_save	[	114	]	;
					tdata_save	[	116	]	<=	tdata_save	[	115	]	;
					tdata_save	[	117	]	<=	tdata_save	[	116	]	;
					tdata_save	[	118	]	<=	tdata_save	[	117	]	;
					tdata_save	[	119	]	<=	tdata_save	[	118	]	;
					tdata_save	[	120	]	<=	tdata_save	[	119	]	;
					tdata_save	[	121	]	<=	tdata_save	[	120	]	;
					tdata_save	[	122	]	<=	tdata_save	[	121	]	;
					tdata_save	[	123	]	<=	tdata_save	[	122	]	;
					tdata_save	[	124	]	<=	tdata_save	[	123	]	;
					tdata_save	[	125	]	<=	tdata_save	[	124	]	;
					tdata_save	[	126	]	<=	tdata_save	[	125	]	;
					tdata_save	[	127	]	<=	tdata_save	[	126	]	;
					tdata_save	[	128	]	<=	tdata_save	[	127	]	;
					tdata_save	[	129	]	<=	tdata_save	[	128	]	;
					tdata_save	[	130	]	<=	tdata_save	[	129	]	;
					tdata_save	[	131	]	<=	tdata_save	[	130	]	;
					tdata_save	[	132	]	<=	tdata_save	[	131	]	;
					tdata_save	[	133	]	<=	tdata_save	[	132	]	;
					tdata_save	[	134	]	<=	tdata_save	[	133	]	;
					tdata_save	[	135	]	<=	tdata_save	[	134	]	;
					tdata_save	[	136	]	<=	tdata_save	[	135	]	;
					tdata_save	[	137	]	<=	tdata_save	[	136	]	;
					tdata_save	[	138	]	<=	tdata_save	[	137	]	;
					tdata_save	[	139	]	<=	tdata_save	[	138	]	;
					tdata_save	[	140	]	<=	tdata_save	[	139	]	;
					tdata_save	[	141	]	<=	tdata_save	[	140	]	;
					tdata_save	[	142	]	<=	tdata_save	[	141	]	;
					tdata_save	[	143	]	<=	tdata_save	[	142	]	;
					tdata_save	[	144	]	<=	tdata_save	[	143	]	;
					tdata_save	[	145	]	<=	tdata_save	[	144	]	;
					tdata_save	[	146	]	<=	tdata_save	[	145	]	;
					tdata_save	[	147	]	<=	tdata_save	[	146	]	;
					tdata_save	[	148	]	<=	tdata_save	[	147	]	;
					tdata_save	[	149	]	<=	tdata_save	[	148	]	;
					tdata_save	[	150	]	<=	tdata_save	[	149	]	;
					tdata_save	[	151	]	<=	tdata_save	[	150	]	;
					tdata_save	[	152	]	<=	tdata_save	[	151	]	;
					tdata_save	[	153	]	<=	tdata_save	[	152	]	;
					tdata_save	[	154	]	<=	tdata_save	[	153	]	;
					tdata_save	[	155	]	<=	tdata_save	[	154	]	;
					tdata_save	[	156	]	<=	tdata_save	[	155	]	;
					tdata_save	[	157	]	<=	tdata_save	[	156	]	;
					tdata_save	[	158	]	<=	tdata_save	[	157	]	;
					tdata_save	[	159	]	<=	tdata_save	[	158	]	;
					tdata_save	[	160	]	<=	tdata_save	[	159	]	;
					tdata_save	[	161	]	<=	tdata_save	[	160	]	;
					tdata_save	[	162	]	<=	tdata_save	[	161	]	;
					tdata_save	[	163	]	<=	tdata_save	[	162	]	;
					tdata_save	[	164	]	<=	tdata_save	[	163	]	;
					tdata_save	[	165	]	<=	tdata_save	[	164	]	;
					tdata_save	[	166	]	<=	tdata_save	[	165	]	;
					tdata_save	[	167	]	<=	tdata_save	[	166	]	;
					tdata_save	[	168	]	<=	tdata_save	[	167	]	;
					tdata_save	[	169	]	<=	tdata_save	[	168	]	;
					tdata_save	[	170	]	<=	tdata_save	[	169	]	;
					tdata_save	[	171	]	<=	tdata_save	[	170	]	;
					tdata_save	[	172	]	<=	tdata_save	[	171	]	;
					tdata_save	[	173	]	<=	tdata_save	[	172	]	;
					tdata_save	[	174	]	<=	tdata_save	[	173	]	;
					tdata_save	[	175	]	<=	tdata_save	[	174	]	;
					tdata_save	[	176	]	<=	tdata_save	[	175	]	;
					tdata_save	[	177	]	<=	tdata_save	[	176	]	;
					tdata_save	[	178	]	<=	tdata_save	[	177	]	;
					tdata_save	[	179	]	<=	tdata_save	[	178	]	;
					tdata_save	[	180	]	<=	tdata_save	[	179	]	;
					tdata_save	[	181	]	<=	tdata_save	[	180	]	;
					tdata_save	[	182	]	<=	tdata_save	[	181	]	;
					tdata_save	[	183	]	<=	tdata_save	[	182	]	;
					tdata_save	[	184	]	<=	tdata_save	[	183	]	;
					tdata_save	[	185	]	<=	tdata_save	[	184	]	;
					tdata_save	[	186	]	<=	tdata_save	[	185	]	;
					tdata_save	[	187	]	<=	tdata_save	[	186	]	;
					tdata_save	[	188	]	<=	tdata_save	[	187	]	;
					tdata_save	[	189	]	<=	tdata_save	[	188	]	;
					tdata_save	[	190	]	<=	tdata_save	[	189	]	;
					tdata_save	[	191	]	<=	tdata_save	[	190	]	;
					tdata_save	[	192	]	<=	tdata_save	[	191	]	;
					tdata_save	[	193	]	<=	tdata_save	[	192	]	;
					tdata_save	[	194	]	<=	tdata_save	[	193	]	;
					tdata_save	[	195	]	<=	tdata_save	[	194	]	;
					tdata_save	[	196	]	<=	tdata_save	[	195	]	;
					tdata_save	[	197	]	<=	tdata_save	[	196	]	;
					tdata_save	[	198	]	<=	tdata_save	[	197	]	;
					tdata_save	[	199	]	<=	tdata_save	[	198	]	;
					tdata_save	[	200	]	<=	tdata_save	[	199	]	;
					tdata_save	[	201	]	<=	tdata_save	[	200	]	;
					tdata_save	[	202	]	<=	tdata_save	[	201	]	;
					tdata_save	[	203	]	<=	tdata_save	[	202	]	;
					tdata_save	[	204	]	<=	tdata_save	[	203	]	;
					tdata_save	[	205	]	<=	tdata_save	[	204	]	;
					tdata_save	[	206	]	<=	tdata_save	[	205	]	;
					tdata_save	[	207	]	<=	tdata_save	[	206	]	;
					tdata_save	[	208	]	<=	tdata_save	[	207	]	;
					tdata_save	[	209	]	<=	tdata_save	[	208	]	;
					tdata_save	[	210	]	<=	tdata_save	[	209	]	;
					tdata_save	[	211	]	<=	tdata_save	[	210	]	;
					tdata_save	[	212	]	<=	tdata_save	[	211	]	;
					tdata_save	[	213	]	<=	tdata_save	[	212	]	;
					tdata_save	[	214	]	<=	tdata_save	[	213	]	;
					tdata_save	[	215	]	<=	tdata_save	[	214	]	;
					tdata_save	[	216	]	<=	tdata_save	[	215	]	;
					tdata_save	[	217	]	<=	tdata_save	[	216	]	;
					tdata_save	[	218	]	<=	tdata_save	[	217	]	;
					tdata_save	[	219	]	<=	tdata_save	[	218	]	;
					tdata_save	[	220	]	<=	tdata_save	[	219	]	;
					tdata_save	[	221	]	<=	tdata_save	[	220	]	;
					tdata_save	[	222	]	<=	tdata_save	[	221	]	;
					tdata_save	[	223	]	<=	tdata_save	[	222	]	;
					tdata_save	[	224	]	<=	tdata_save	[	223	]	;
					tdata_save	[	225	]	<=	tdata_save	[	224	]	;
					tdata_save	[	226	]	<=	tdata_save	[	225	]	;
					tdata_save	[	227	]	<=	tdata_save	[	226	]	;
					tdata_save	[	228	]	<=	tdata_save	[	227	]	;
					tdata_save	[	229	]	<=	tdata_save	[	228	]	;
					tdata_save	[	230	]	<=	tdata_save	[	229	]	;
					tdata_save	[	231	]	<=	tdata_save	[	230	]	;
					tdata_save	[	232	]	<=	tdata_save	[	231	]	;
					tdata_save	[	233	]	<=	tdata_save	[	232	]	;
					tdata_save	[	234	]	<=	tdata_save	[	233	]	;
					tdata_save	[	235	]	<=	tdata_save	[	234	]	;
					tdata_save	[	236	]	<=	tdata_save	[	235	]	;
					tdata_save	[	237	]	<=	tdata_save	[	236	]	;
					tdata_save	[	238	]	<=	tdata_save	[	237	]	;
					tdata_save	[	239	]	<=	tdata_save	[	238	]	;
					tdata_save	[	240	]	<=	tdata_save	[	239	]	;
					tdata_save	[	241	]	<=	tdata_save	[	240	]	;
					tdata_save	[	242	]	<=	tdata_save	[	241	]	;
					tdata_save	[	243	]	<=	tdata_save	[	242	]	;
					tdata_save	[	244	]	<=	tdata_save	[	243	]	;
					tdata_save	[	245	]	<=	tdata_save	[	244	]	;
					tdata_save	[	246	]	<=	tdata_save	[	245	]	;
					tdata_save	[	247	]	<=	tdata_save	[	246	]	;
					tdata_save	[	248	]	<=	tdata_save	[	247	]	;
					tdata_save	[	249	]	<=	tdata_save	[	248	]	;
					tdata_save	[	250	]	<=	tdata_save	[	249	]	;
					tdata_save	[	251	]	<=	tdata_save	[	250	]	;
					tdata_save	[	252	]	<=	tdata_save	[	251	]	;
					tdata_save	[	253	]	<=	tdata_save	[	252	]	;
					tdata_save	[	254	]	<=	tdata_save	[	253	]	;
					tdata_save	[	255	]	<=	tdata_save	[	254	]	;
					tuser_save	[	0	]	<=	tuser;						
				tuser_save	[	1	]	<=	tuser_save	[	0	]	;
				tuser_save	[	2	]	<=	tuser_save	[	1	]	;
				tuser_save	[	3	]	<=	tuser_save	[	2	]	;
				tuser_save	[	4	]	<=	tuser_save	[	3	]	;
				tuser_save	[	5	]	<=	tuser_save	[	4	]	;
				tuser_save	[	6	]	<=	tuser_save	[	5	]	;
				tuser_save	[	7	]	<=	tuser_save	[	6	]	;
				tuser_save	[	8	]	<=	tuser_save	[	7	]	;
				tuser_save	[	9	]	<=	tuser_save	[	8	]	;
				tuser_save	[	10	]	<=	tuser_save	[	9	]	;
				tuser_save	[	11	]	<=	tuser_save	[	10	]	;
				tuser_save	[	12	]	<=	tuser_save	[	11	]	;
				tuser_save	[	13	]	<=	tuser_save	[	12	]	;
				tuser_save	[	14	]	<=	tuser_save	[	13	]	;
				tuser_save	[	15	]	<=	tuser_save	[	14	]	;
				tuser_save	[	16	]	<=	tuser_save	[	15	]	;
				tuser_save	[	17	]	<=	tuser_save	[	16	]	;
				tuser_save	[	18	]	<=	tuser_save	[	17	]	;
				tuser_save	[	19	]	<=	tuser_save	[	18	]	;
				tuser_save	[	20	]	<=	tuser_save	[	19	]	;
				tuser_save	[	21	]	<=	tuser_save	[	20	]	;
				tuser_save	[	22	]	<=	tuser_save	[	21	]	;
				tuser_save	[	23	]	<=	tuser_save	[	22	]	;
				tuser_save	[	24	]	<=	tuser_save	[	23	]	;
				tuser_save	[	25	]	<=	tuser_save	[	24	]	;
				tuser_save	[	26	]	<=	tuser_save	[	25	]	;
				tuser_save	[	27	]	<=	tuser_save	[	26	]	;
				tuser_save	[	28	]	<=	tuser_save	[	27	]	;
				tuser_save	[	29	]	<=	tuser_save	[	28	]	;
				tuser_save	[	30	]	<=	tuser_save	[	29	]	;
				tuser_save	[	31	]	<=	tuser_save	[	30	]	;
				tuser_save	[	32	]	<=	tuser_save	[	31	]	;
				tuser_save	[	33	]	<=	tuser_save	[	32	]	;
				tuser_save	[	34	]	<=	tuser_save	[	33	]	;
				tuser_save	[	35	]	<=	tuser_save	[	34	]	;
				tuser_save	[	36	]	<=	tuser_save	[	35	]	;
				tuser_save	[	37	]	<=	tuser_save	[	36	]	;
				tuser_save	[	38	]	<=	tuser_save	[	37	]	;
				tuser_save	[	39	]	<=	tuser_save	[	38	]	;
				tuser_save	[	40	]	<=	tuser_save	[	39	]	;
				tuser_save	[	41	]	<=	tuser_save	[	40	]	;
				tuser_save	[	42	]	<=	tuser_save	[	41	]	;
				tuser_save	[	43	]	<=	tuser_save	[	42	]	;
				tuser_save	[	44	]	<=	tuser_save	[	43	]	;
				tuser_save	[	45	]	<=	tuser_save	[	44	]	;
				tuser_save	[	46	]	<=	tuser_save	[	45	]	;
				tuser_save	[	47	]	<=	tuser_save	[	46	]	;
				tuser_save	[	48	]	<=	tuser_save	[	47	]	;
				tuser_save	[	49	]	<=	tuser_save	[	48	]	;
				tuser_save	[	50	]	<=	tuser_save	[	49	]	;
				tuser_save	[	51	]	<=	tuser_save	[	50	]	;
				tuser_save	[	52	]	<=	tuser_save	[	51	]	;
				tuser_save	[	53	]	<=	tuser_save	[	52	]	;
				tuser_save	[	54	]	<=	tuser_save	[	53	]	;
				tuser_save	[	55	]	<=	tuser_save	[	54	]	;
				tuser_save	[	56	]	<=	tuser_save	[	55	]	;
				tuser_save	[	57	]	<=	tuser_save	[	56	]	;
				tuser_save	[	58	]	<=	tuser_save	[	57	]	;
				tuser_save	[	59	]	<=	tuser_save	[	58	]	;
				tuser_save	[	60	]	<=	tuser_save	[	59	]	;
				tuser_save	[	61	]	<=	tuser_save	[	60	]	;
				tuser_save	[	62	]	<=	tuser_save	[	61	]	;
				tuser_save	[	63	]	<=	tuser_save	[	62	]	;
				tuser_save	[	64	]	<=	tuser_save	[	63	]	;
				tuser_save	[	65	]	<=	tuser_save	[	64	]	;
				tuser_save	[	66	]	<=	tuser_save	[	65	]	;
				tuser_save	[	67	]	<=	tuser_save	[	66	]	;
				tuser_save	[	68	]	<=	tuser_save	[	67	]	;
				tuser_save	[	69	]	<=	tuser_save	[	68	]	;
				tuser_save	[	70	]	<=	tuser_save	[	69	]	;
				tuser_save	[	71	]	<=	tuser_save	[	70	]	;
				tuser_save	[	72	]	<=	tuser_save	[	71	]	;
				tuser_save	[	73	]	<=	tuser_save	[	72	]	;
				tuser_save	[	74	]	<=	tuser_save	[	73	]	;
				tuser_save	[	75	]	<=	tuser_save	[	74	]	;
				tuser_save	[	76	]	<=	tuser_save	[	75	]	;
				tuser_save	[	77	]	<=	tuser_save	[	76	]	;
				tuser_save	[	78	]	<=	tuser_save	[	77	]	;
				tuser_save	[	79	]	<=	tuser_save	[	78	]	;
				tuser_save	[	80	]	<=	tuser_save	[	79	]	;
				tuser_save	[	81	]	<=	tuser_save	[	80	]	;
				tuser_save	[	82	]	<=	tuser_save	[	81	]	;
				tuser_save	[	83	]	<=	tuser_save	[	82	]	;
				tuser_save	[	84	]	<=	tuser_save	[	83	]	;
				tuser_save	[	85	]	<=	tuser_save	[	84	]	;
				tuser_save	[	86	]	<=	tuser_save	[	85	]	;
				tuser_save	[	87	]	<=	tuser_save	[	86	]	;
				tuser_save	[	88	]	<=	tuser_save	[	87	]	;
				tuser_save	[	89	]	<=	tuser_save	[	88	]	;
				tuser_save	[	90	]	<=	tuser_save	[	89	]	;
				tuser_save	[	91	]	<=	tuser_save	[	90	]	;
				tuser_save	[	92	]	<=	tuser_save	[	91	]	;
				tuser_save	[	93	]	<=	tuser_save	[	92	]	;
				tuser_save	[	94	]	<=	tuser_save	[	93	]	;
				tuser_save	[	95	]	<=	tuser_save	[	94	]	;
				tuser_save	[	96	]	<=	tuser_save	[	95	]	;
				tuser_save	[	97	]	<=	tuser_save	[	96	]	;
				tuser_save	[	98	]	<=	tuser_save	[	97	]	;
				tuser_save	[	99	]	<=	tuser_save	[	98	]	;
				tuser_save	[	100	]	<=	tuser_save	[	99	]	;
				tuser_save	[	101	]	<=	tuser_save	[	100	]	;
				tuser_save	[	102	]	<=	tuser_save	[	101	]	;
				tuser_save	[	103	]	<=	tuser_save	[	102	]	;
				tuser_save	[	104	]	<=	tuser_save	[	103	]	;
				tuser_save	[	105	]	<=	tuser_save	[	104	]	;
				tuser_save	[	106	]	<=	tuser_save	[	105	]	;
				tuser_save	[	107	]	<=	tuser_save	[	106	]	;
				tuser_save	[	108	]	<=	tuser_save	[	107	]	;
				tuser_save	[	109	]	<=	tuser_save	[	108	]	;
				tuser_save	[	110	]	<=	tuser_save	[	109	]	;
				tuser_save	[	111	]	<=	tuser_save	[	110	]	;
				tuser_save	[	112	]	<=	tuser_save	[	111	]	;
				tuser_save	[	113	]	<=	tuser_save	[	112	]	;
				tuser_save	[	114	]	<=	tuser_save	[	113	]	;
				tuser_save	[	115	]	<=	tuser_save	[	114	]	;
				tuser_save	[	116	]	<=	tuser_save	[	115	]	;
				tuser_save	[	117	]	<=	tuser_save	[	116	]	;
				tuser_save	[	118	]	<=	tuser_save	[	117	]	;
				tuser_save	[	119	]	<=	tuser_save	[	118	]	;
				tuser_save	[	120	]	<=	tuser_save	[	119	]	;
				tuser_save	[	121	]	<=	tuser_save	[	120	]	;
				tuser_save	[	122	]	<=	tuser_save	[	121	]	;
				tuser_save	[	123	]	<=	tuser_save	[	122	]	;
				tuser_save	[	124	]	<=	tuser_save	[	123	]	;
				tuser_save	[	125	]	<=	tuser_save	[	124	]	;
				tuser_save	[	126	]	<=	tuser_save	[	125	]	;
				tuser_save	[	127	]	<=	tuser_save	[	126	]	;
				tuser_save	[	128	]	<=	tuser_save	[	127	]	;
				tuser_save	[	129	]	<=	tuser_save	[	128	]	;
				tuser_save	[	130	]	<=	tuser_save	[	129	]	;
				tuser_save	[	131	]	<=	tuser_save	[	130	]	;
				tuser_save	[	132	]	<=	tuser_save	[	131	]	;
				tuser_save	[	133	]	<=	tuser_save	[	132	]	;
				tuser_save	[	134	]	<=	tuser_save	[	133	]	;
				tuser_save	[	135	]	<=	tuser_save	[	134	]	;
				tuser_save	[	136	]	<=	tuser_save	[	135	]	;
				tuser_save	[	137	]	<=	tuser_save	[	136	]	;
				tuser_save	[	138	]	<=	tuser_save	[	137	]	;
				tuser_save	[	139	]	<=	tuser_save	[	138	]	;
				tuser_save	[	140	]	<=	tuser_save	[	139	]	;
				tuser_save	[	141	]	<=	tuser_save	[	140	]	;
				tuser_save	[	142	]	<=	tuser_save	[	141	]	;
				tuser_save	[	143	]	<=	tuser_save	[	142	]	;
				tuser_save	[	144	]	<=	tuser_save	[	143	]	;
				tuser_save	[	145	]	<=	tuser_save	[	144	]	;
				tuser_save	[	146	]	<=	tuser_save	[	145	]	;
				tuser_save	[	147	]	<=	tuser_save	[	146	]	;
				tuser_save	[	148	]	<=	tuser_save	[	147	]	;
				tuser_save	[	149	]	<=	tuser_save	[	148	]	;
				tuser_save	[	150	]	<=	tuser_save	[	149	]	;
				tuser_save	[	151	]	<=	tuser_save	[	150	]	;
				tuser_save	[	152	]	<=	tuser_save	[	151	]	;
				tuser_save	[	153	]	<=	tuser_save	[	152	]	;
				tuser_save	[	154	]	<=	tuser_save	[	153	]	;
				tuser_save	[	155	]	<=	tuser_save	[	154	]	;
				tuser_save	[	156	]	<=	tuser_save	[	155	]	;
				tuser_save	[	157	]	<=	tuser_save	[	156	]	;
				tuser_save	[	158	]	<=	tuser_save	[	157	]	;
				tuser_save	[	159	]	<=	tuser_save	[	158	]	;
				tuser_save	[	160	]	<=	tuser_save	[	159	]	;
				tuser_save	[	161	]	<=	tuser_save	[	160	]	;
				tuser_save	[	162	]	<=	tuser_save	[	161	]	;
				tuser_save	[	163	]	<=	tuser_save	[	162	]	;
				tuser_save	[	164	]	<=	tuser_save	[	163	]	;
				tuser_save	[	165	]	<=	tuser_save	[	164	]	;
				tuser_save	[	166	]	<=	tuser_save	[	165	]	;
				tuser_save	[	167	]	<=	tuser_save	[	166	]	;
				tuser_save	[	168	]	<=	tuser_save	[	167	]	;
				tuser_save	[	169	]	<=	tuser_save	[	168	]	;
				tuser_save	[	170	]	<=	tuser_save	[	169	]	;
				tuser_save	[	171	]	<=	tuser_save	[	170	]	;
				tuser_save	[	172	]	<=	tuser_save	[	171	]	;
				tuser_save	[	173	]	<=	tuser_save	[	172	]	;
				tuser_save	[	174	]	<=	tuser_save	[	173	]	;
				tuser_save	[	175	]	<=	tuser_save	[	174	]	;
				tuser_save	[	176	]	<=	tuser_save	[	175	]	;
				tuser_save	[	177	]	<=	tuser_save	[	176	]	;
				tuser_save	[	178	]	<=	tuser_save	[	177	]	;
				tuser_save	[	179	]	<=	tuser_save	[	178	]	;
				tuser_save	[	180	]	<=	tuser_save	[	179	]	;
				tuser_save	[	181	]	<=	tuser_save	[	180	]	;
				tuser_save	[	182	]	<=	tuser_save	[	181	]	;
				tuser_save	[	183	]	<=	tuser_save	[	182	]	;
				tuser_save	[	184	]	<=	tuser_save	[	183	]	;
				tuser_save	[	185	]	<=	tuser_save	[	184	]	;
				tuser_save	[	186	]	<=	tuser_save	[	185	]	;
				tuser_save	[	187	]	<=	tuser_save	[	186	]	;
				tuser_save	[	188	]	<=	tuser_save	[	187	]	;
				tuser_save	[	189	]	<=	tuser_save	[	188	]	;
				tuser_save	[	190	]	<=	tuser_save	[	189	]	;
				tuser_save	[	191	]	<=	tuser_save	[	190	]	;
				tuser_save	[	192	]	<=	tuser_save	[	191	]	;
				tuser_save	[	193	]	<=	tuser_save	[	192	]	;
				tuser_save	[	194	]	<=	tuser_save	[	193	]	;
				tuser_save	[	195	]	<=	tuser_save	[	194	]	;
				tuser_save	[	196	]	<=	tuser_save	[	195	]	;
				tuser_save	[	197	]	<=	tuser_save	[	196	]	;
				tuser_save	[	198	]	<=	tuser_save	[	197	]	;
				tuser_save	[	199	]	<=	tuser_save	[	198	]	;
				tuser_save	[	200	]	<=	tuser_save	[	199	]	;
				tuser_save	[	201	]	<=	tuser_save	[	200	]	;
				tuser_save	[	202	]	<=	tuser_save	[	201	]	;
				tuser_save	[	203	]	<=	tuser_save	[	202	]	;
				tuser_save	[	204	]	<=	tuser_save	[	203	]	;
				tuser_save	[	205	]	<=	tuser_save	[	204	]	;
				tuser_save	[	206	]	<=	tuser_save	[	205	]	;
				tuser_save	[	207	]	<=	tuser_save	[	206	]	;
				tuser_save	[	208	]	<=	tuser_save	[	207	]	;
				tuser_save	[	209	]	<=	tuser_save	[	208	]	;
				tuser_save	[	210	]	<=	tuser_save	[	209	]	;
				tuser_save	[	211	]	<=	tuser_save	[	210	]	;
				tuser_save	[	212	]	<=	tuser_save	[	211	]	;
				tuser_save	[	213	]	<=	tuser_save	[	212	]	;
				tuser_save	[	214	]	<=	tuser_save	[	213	]	;
				tuser_save	[	215	]	<=	tuser_save	[	214	]	;
				tuser_save	[	216	]	<=	tuser_save	[	215	]	;
				tuser_save	[	217	]	<=	tuser_save	[	216	]	;
				tuser_save	[	218	]	<=	tuser_save	[	217	]	;
				tuser_save	[	219	]	<=	tuser_save	[	218	]	;
				tuser_save	[	220	]	<=	tuser_save	[	219	]	;
				tuser_save	[	221	]	<=	tuser_save	[	220	]	;
				tuser_save	[	222	]	<=	tuser_save	[	221	]	;
				tuser_save	[	223	]	<=	tuser_save	[	222	]	;
				tuser_save	[	224	]	<=	tuser_save	[	223	]	;
				tuser_save	[	225	]	<=	tuser_save	[	224	]	;
				tuser_save	[	226	]	<=	tuser_save	[	225	]	;
				tuser_save	[	227	]	<=	tuser_save	[	226	]	;
				tuser_save	[	228	]	<=	tuser_save	[	227	]	;
				tuser_save	[	229	]	<=	tuser_save	[	228	]	;
				tuser_save	[	230	]	<=	tuser_save	[	229	]	;
				tuser_save	[	231	]	<=	tuser_save	[	230	]	;
				tuser_save	[	232	]	<=	tuser_save	[	231	]	;
				tuser_save	[	233	]	<=	tuser_save	[	232	]	;
				tuser_save	[	234	]	<=	tuser_save	[	233	]	;
				tuser_save	[	235	]	<=	tuser_save	[	234	]	;
				tuser_save	[	236	]	<=	tuser_save	[	235	]	;
				tuser_save	[	237	]	<=	tuser_save	[	236	]	;
				tuser_save	[	238	]	<=	tuser_save	[	237	]	;
				tuser_save	[	239	]	<=	tuser_save	[	238	]	;
				tuser_save	[	240	]	<=	tuser_save	[	239	]	;
				tuser_save	[	241	]	<=	tuser_save	[	240	]	;
				tuser_save	[	242	]	<=	tuser_save	[	241	]	;
				tuser_save	[	243	]	<=	tuser_save	[	242	]	;
				tuser_save	[	244	]	<=	tuser_save	[	243	]	;
				tuser_save	[	245	]	<=	tuser_save	[	244	]	;
				tuser_save	[	246	]	<=	tuser_save	[	245	]	;
				tuser_save	[	247	]	<=	tuser_save	[	246	]	;
				tuser_save	[	248	]	<=	tuser_save	[	247	]	;
				tuser_save	[	249	]	<=	tuser_save	[	248	]	;
				tuser_save	[	250	]	<=	tuser_save	[	249	]	;
				tuser_save	[	251	]	<=	tuser_save	[	250	]	;
				tuser_save	[	252	]	<=	tuser_save	[	251	]	;
				tuser_save	[	253	]	<=	tuser_save	[	252	]	;
				tuser_save	[	254	]	<=	tuser_save	[	253	]	;
				tuser_save	[	255	]	<=	tuser_save	[	254	]	;
				if(count_packet == 2'd2)
				begin
					count_packet <= 2'd0;
				end
				else
				begin
					count_packet	<= count_packet;
				end
				sum_tdata		<=	tdata_save[255];
				sum_tuser		<=	tuser_save[127];
				sum_tdata_valid		<=	1'b1;
				sum_tuser_valid		<=	1'b1;
			end
		end
	end
		
	//axi to fifo --> asyc_fifo read enable
	always@(*)
	begin
		inc = axififo_din_valid && ((~axififo_empty) && ~axififo_mem_queue_full);
		inc_tuser = dout_valid_tuser && ((~rempty_tuser) && ~axififo_mem_queue_full);
	end

endmodule

